`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JuD9eDvwcSlj3mddIdgx2eU7vtHTUReS3Iu5T4oCZYwRlea8s4rn8AGQ7Z7jxB+zHF93LIe3s+ZK
1PT7VHtdNQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B6MSz4lAKwGigp7QQp9aE8dHAFnYn+aoNN5DtGimC7WTUCQhHIdvVo1byuDtfzlmGCM6OuyKuPpS
8cONvqFyv51r7L+amtJ+UgplwqG1EDv4HHx4XZuHypuor2F5DRZ8I3La36ehF4fr6cnJdnoB9ofv
yNMx3aNvdjXtKIGL4Uk=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Gr1L/7sTpu+m3XYWbedbgoUJkl3VdNRB+c23FmidnFV2lEukogbcs3BbUuKAV/PQh3jaB+51lm5E
Wpl+dpv3FqgytzDwLS/ClSU7xwgc49nLV6gUYMZ+IwfPVp4p17iuhK4NFPPnNHdHpq9bpRJ7i7qv
23zVJxXmmF1Hb7n9B1N3KHDCgPF4z3UDXb690K0IaXwji9FjYNgW+Zu1HKm3kQJMoSw0D38q0tDb
WKtE8dDselx/BlaodG7RpHiAFDQmWwgNGQyWK8iy2HHaaGUR0rxqM/dqtcviAIiXB9QNnPG/Kow1
udoLyxpr9OnpTj9Eotttc0uF0bW13Zq2OL7Skg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u4sdiAb6lY4dwm5aYaJzX4XbGcLIYsX5R9yeM7SvtO4l/gsdRnn+bAXWg36RhrG1v3G3hfQJt+Re
uUsRONch5aWmR0XXVof+Ak7T8Sbb4k5zrLuO4Nl0vu/vP2TyQDYSYvPpkYZfb0wcdZJcH3trN6TZ
hd1XdPBnwBIAigqolmTdSmsRynoqmc73oJbJMlIn792oevR2RL2eqM5q/9UgC4CC45Avk4fTpXPn
0c5AeOkKiwxawRbJE8qCro2DrgE4NKePwHqh36a2Hvv/JfyF30D/PBeX5/NMhjZoHCkIFthBU3p/
NDpXoe1prXrQjgFSpi7xpkiC0eiS9ZZyCls5sA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Xf9IdAuk+kSAJlBFFF2Aqc4wHLr8efsHLyp/13z6rPpqorq0OfQDApTV9XSKi7DMMN88Ny+Rrb2j
5amLfWsqfH8DASPGGVuWp5K+CDGbLCCvfotVpwfvlcwCKHAMsTn4FXcq2JSIHGhNr2NiF0s9GjFV
63wTuCBpnbG0qmdAL239JN90hu424LUSg93v94XQA+PRHNpgRWZclIo1fggKtO0uveTdo5Q6/7Vb
b1kU+p8xUQhnzUuNnZ/b5uG/hiCbiEUsbaXnOv7DY6/Qbn1BjlKtyC4hPUeLxPkH/6VvdwyV7Y+f
KuaJ8GZ3JWRgMX22rF9S+CNsiNfnkDhJprWWDA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ia3x9ja6nx2nE1syG5TIYkxEErHOHGaJgnLU9baMpfhOT+/Nq64lrSsmvf/0dNJOpqrV/CO3Jhox
0f8JYxWbrUSksd98ku2xyZOpk0MsBiPYM89NTIIA1+CXJbkpGGnel9Wz3WHr8Xu3YeydDeymqoc6
IXJLFFYa5Rzjn+ls6qo=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LJwNWX8uWfXzsQK1ukh51ZJbvpWFk0mZuuoxfOh2NbOhgFmIt6b06CkJtFYygrc/ZXI3LgwHQUWp
A3XxGmUMnGrEiFBTMXHll3ViO/Jj5vd/uQue0q8UwMLCwNcafOShfIqeMhfDvbk+s8SBiXFmply4
MWBZ1YbL8faiFb8WVWSDkchm4TekKbKdeqzu8H0mj+PBhE4VNJJnBvNlplcSkT1JoW99HTxln8u5
aV/n66LZRmoPMSNpR30HL4FC8eaUDAQutAIR9nGSJRJFuU7jHih0x0ixgW2Wx4/D1MU1haxZM1u/
dxzNlK7OREy7OswIfsbxFxbmIqywf4CFk10QJA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57632)
`protect data_block
DaJymrSD1FYBFG7UVcmZkm2iYVYImxJz1/u5245JOOOzBaxz0QlGZaWg+2YsnGg9k6wP3L8iMi0s
k1xhPuqCZB8MXz/zhjQbfwEnq5ES9P6hEV9xyU0hqre0NXWfY5iNgmJ+spCKVlRJ7EULm8bsA9QH
8SFOYBHDBugIsb1z994NteZRiJCtQ2dCVA8IQxyxtth7elYwfVIxHeW23XNcTXowpC79C0QqfV82
nati8C1id4VkJeaEfslYEQ0wEu7nx6iAXAW3vd8nFLC/84a3dn0ngG1l9CfDXrU+rSYay75fDfNZ
gQSRYM2C0ui/YSztJZC8dKaWNKiGnkClnm77exYSrTFkdJKzGnNv6kM7SZipXmYViVrp36VSkzyb
LZppO730Zg1JZi6bOv3zEoaBuGgOKY29IS5RGbVeDBgd+gHoNW3fdKGoyIZ8WZ+bivFnD4p1OFnr
R3NvoS181wFNiNAIdycDEk8abDj8MEH+drWapIrr3B0TO5y28bbOjsUiEQWXjE8XDl6f6Di9Rjag
uPoScNjJXSXPeu15MDPdCKDzYYPH8VAHpJfBfXi11mtNCZ7PytyrskvbW7mZA+vbrc1d+jUy/T3f
MBGkhHFKBPlsSiASxVZDe1pcCb7isZQVOAN3N5wjMldSE9MMahHUiiXNWkoCHnK4yTItz19j8zEz
G4XPhjmkthtfuZ04Odf3t0ic8aWVQUvVGd5IVaJOUEk1DvfHqmxuGijF1fVJJNDXC0MYDvRJzJ6z
3ZVhq+qOqevYXMfxOWd5kgAAQ6Qlr9Sw/+INiYHIY3oD46kB6dt2jAvnmePlux9VnXwBDkC+uOsK
9b6Hzas7RrxW6MUR7x9dUXW/QfdnFSzlCI9NUynbrvWByu06iaFa8zyRD4tZitX+2DdUl7c+8tPX
KJEF4aei7GgP/yP4hkqiqK2teLaCicMoe/eTwCp/aWL3hGwKlks79B0qfdMI3T3echX7NY8cv23x
ejwxBiZ/CTAAOVJRW9ObbABtdFZPQiZ1xkejglEnsLZYkWY/F49X5CGuux4FdKfgRmEK1qCHyzU8
EaR7zAmnyGnlee7qdls9jCVZmadDvfvEAARMD9Bj+YNmXcAgjj6JKC6iwtD52TpOwtscMXXqlN0H
dxx49YHdES3KP+gMkPaKQz2uQgDacyHbW5CmjyzcmR0SFQYAwbCEFNjkmhlrEfVLFo0so/fOmYZl
uJxmF3KVzW26aKQdyXN3299J1sNmIfx0t2WCLwquK097d+aowk5R94LiMZnMP9Yj54ANPk2W17uM
H6LdKSQL3L7AfePcQuZF3SCycO6RVqk43TcKqdDU1AH6mt643FIRleF4ZwBL7tkSUM2l4HTcnVtN
mlbbSDKVj+zjBw/VJIX3C4oda/hyJm9aB3AIttcXBWFMR3urwoRTdimgcOawM7TproMTzsbkdCk4
l2P+hOF/vzevmZ+R7td097pBVLUMt0t1uhMy3N9kG0t10V/d4PwjfG2trFJKlt9nyV4gCuVhBwjI
86M+MyrIVFcvB1DWBQX9TE8+okQ/X+e5ra81o2P/DwZGFbYj5Vd3DR8yDyRQoHAws+w9m6T81d4h
pfAZNHcqB0pstgFMdyQEh0E5UTXhItgC/0CSpeYRbXatZNMm033Tj/R/sw0YnQh8P2J/oEMokIGq
ngJwQ9hUpAUhriPewYEfxW0+2x97K7geXMwxGtEXUolncX3AVrt4vhE7NH4eLcto1eCT+IGoKLAZ
j3z+CFbWQFgHquQ2aHfA3C7O6FbTqDNzhrnF400IMo/muhLBHN9yfTlLulo8bQBs/xMl4quwgeqO
LeaQiZZ9F0uMgujYzrTmMnzao6oqFgnz6C5v+wbYqOBCgDzMkOg55PuRUSmbRAJ+NbOkPK1rzePi
oM4Phygvd6ahNXYk4uF4hYz2ZcypLXdv4Oa2QIkZxmwrPtWQQ9BO3fxn6UgDqSWX+NmZPTLzClWb
qrOWu3EJU+mxjrYDq1F/hqrEcHF8XjqC3diVXfk1PViT3ChkCPzhRVCzMekvbVzo649awbwjqnSR
Gx9PdIA5mmzyMIHsKr+zj0NaCuu3XoDAOLm9FN/GV71Dyz2cavwbCeqTku9ylK5DdxsYhz2jYTHh
0h6ZXKXks5+SKEUYavRzFTlLIiwQckxZLrJiv0mlTeOD2vci2vB3sBJc/XJ+HJeKTD4CH5vg0MEU
deYqlRMK/elvTkadJGYrIH7RIK06Is9DN1qdWqQTu9S3Ll3Len/0fzwJ5UhYbMid8CYAu0aGuAjJ
OuNFyQtHlL/hSOQavCGj8GUZ2u1cB9d9dk9F88ZvC9JBfDNAMMIKblP6mEz5Ke/bHyBH577oHLMf
sjzRJvEwV3I5fEtJyDxsGRkWv8ZM38wQCBSMIDFsZ7owAkaJ8HVzQuQYKhegZ54YX7k9PCvWpKJr
Fa/IAFtjKIvB0DNKrQnji4+LsIhLgd0fKYZDpYzQl2n4GFkj6oc9/fpR8qEObFhdsuaXrkjRh43C
jPAKQOP5dKHDzD3ApK3bRqCyb2G/F8eZCa35xKxPgje6TKffVJzG5AA7Zhs1zplvxztguxWnji87
wI5TYWAON1BSwgLhMExfOeNZt49T2EYMFOWUB5OUjXm3tEtHZkNPQviCYj85luqInoBhEYCH7opj
A56qWQPR8i4CNzHOVgb/6s6nYsP0u8fxVgAUO7ZUamdzaIIgHSz8uVWc0W8sgbzEC3alGqycU4lo
rPkUgCwJoiydOHP+D2scnCM3+U5ylvQS3eZ4Pdm2hMNbeaOEaKcLzY5m1aIIlRNcCUqim1TAymMe
dPknr0r6emtZxAaEJf2J2dsQFrktaIH7YRu15jutYM6wZaTGBlsg16RHKqAcQiZRB+d/HzybzHIU
F3ktvwRvtQvDhhpg0HKXDwBgmFliELvpu0io+w1+LW3mrhwwpx7S4mB+my0n8qCB8iI24z3Qalwn
tf4gx3mGiNAKGgxGFYtbZo9K1qXj+OXVULmm+oEhuLFIimRN3sS3jz6ZK/LUPIAYuI7wkfwRc+d4
G2fLgcRvYgssO5N2yDGg7mK/aQaKGI+mmjmG38pOGaE9R3qHyJ8cnynd2JZMPP8PQ/yBBe9OfTNE
zpNyg1KAutVJ+8lANYJr5Vbx7aAURzpm9Ci7kVM8sk4D61FtZBVh8YfLCYM57jUBmUOi6ZICbouh
jZfV/2mO+GpmdHdb7qUgU7CVTGDBLm7M/JXX6NX1hVXc0eFAZJnUrqsGTcgiq9Sa/iKpbh3GN5gh
KN6JdPFy5kTcctv2gnWNiQSZvW+RDc59mwM7EuYQfNUltlqvYjDYEGXmoaMCBfyHIC3370xavY8E
qR2/xwJH2bjvU+Dwr7Jl40/L3ZIDMKKEqSfHm0r1x48+LcWM3aK9DQ7EJ0n2s5IY31b/s4C8dsns
X9FwSWrWcIkmdSbNm56tBuksZ2fD3r08zLmaB5T5bCvAv/si43jy4PtL/WbiQsMu6W9BnB2CXamL
NnEsp+UhK1ahimgUoK8SjXBVphWUpxMblvmJFTRA+OBAKAB3iRVRcnDj+KuutQaH3SbBB7qcd+JD
PUVNSuFDGUQi4DXigJmgGw5QkEFEH8jAsCfo1efdNJmKzvfiBu9o6L91eSLMKIZ8XUGh64dyQj7p
6Qvv9YhdOzy1eOMKuCj/COmzNI6bDNKARWUEJmmiD7He5zepgrT+KHprt4+IRMlHSlc1RSk4czJP
4fkSYOrbMMVdzNIGzBOeKNg4UCOejt+4PayoQd60Hr8ae1eNaWaTfz3pMx9ZF1QK/+7PtOcg5LiI
2/lnoj5gmG5U1ANcoi+idAqivc/r5At0dwLL5UBw4FzuMeEDBO0r4SD2dTUvim68Sk2HESXOWIQA
RL+VA52mF6lg5EYSlVe7PUykGrY4moV+mq8mQ7RHBE9dweDKJ4QB8C/c/nTf+Y/5SIPvbtG1Str7
KR0dWPcQDDkVzqAra9MgAHxm4x63QYwXCa5vgpI1cY13gRvd6ZbzYZr2ZGbgFfgD/FHr6zgQMYRq
3GGmzQLT+nx19Aw05w1R0Dajmq86r609BAPD9R8IzYDrB3NvHSuuT3KRrq9koVkkEXHewsCbNF0v
h6WxrJwBEYVOcm8YumsTEtAJq5/iJZSaroGQ9ZtGCkCgu0cYYFrX9zJ9vF79ZN2MDJYqW6f/iZ9T
H5PC6ErMMsZ3SWe1+Xoq2qC1VdrMQS8lCplIfHgb7c/ljXaXU68NQQ66seHYx4Ox3zEPcEmnl45o
ZOGzPrmE8RgfR5stxqNJxu0arCOsP+EVkzMCH3cIUvQi7g7bQ7KGQcMU28X/cmEv+vxKopaW4Evy
w+KHjfzTPo8fFglUerqDxeARUSIiFW5GmjcBw1ycBYe4vV+WHOi/hUjspuysvRZX2UTjtiuPyybl
GpgMKyBW8N2BViytDK2X9MceoWVjssAbSdSXUCqYnNY6XDTQkPVtsP4JS6VIrOiF6h08vpPORb6i
FUVOuC1wf26FrLJb79SBiMvu/R//ZwN6Og2s2Dl393cnIu/Uo1Rbj79Pd4Y5bjq0Ufx6N5so4HBL
aNP1+Y3h+yBN06BucJ5G1Gk69SpMEiQ0Fd84IaQesLRhzEsriHQBfVJHe603LbwBQytpUxCUO+WM
f/mwPDdvCkkGUk1REpIivqwNz17KuGrnmHOZUvEOSDE0+BrvysTVhqEnxy4PEwnM8cWKWItBD/ek
tCTeZpQ2wsqNV80axgvfel1NGaarpvV9zEbS4FNI1sDWHQfDQe1jWCDNdDog9OjnRtaTdEr1WW3w
bSOPoUh0M+SQZhx+MtD0sg05Zb6LSu6t3sGJWXpY9qjvzHvlBJ7HqApQOFW0F9P6bJ4gKR1uQ/U3
b0+Mws21IzRN6RI1q/3PVOcAv7eRtPqCpT7Radp8bjRZvR3DTKMSCi8KGkrbesgF83bCehmec38W
LSww1swl4n09DZrHJsWFtwNeStd5LXwr6qVLCsG4dXjkVm6AdwgvUPGbQqtsC316z3CSwGlVJT/t
LaGBti/9GTnpn01q1Yed7fd5vpHLUHl5poLDREq73vCUyRK33Fw4iP7iny/L2EeEar8NcYGl/2TQ
mzkWFw0k1JpRn+85eWPRROCUBAxs41N8fRcrfST0Yp2J1lXM7gcJbnW/dm3wDDhNhg6QeKgiqETi
JbdlcEkHlUWV5qYHNb5u67BifDpWY/PPoZoYtIi5EYGhdsJ0pHv7OvNe3cm8KftwVI9eKsQXuAn+
4UUGx/yWuhl5LWw3z264Ma/hwvjIqX310hR3blYCjHLOpaCqIoFpwCTSzdXAz4h2NTpLuDMG94Zf
sguTWPMvCJZthAw2r7y84rZzSBwEwUStmaYSHS5nZMJr9qMuO7LQivUT1I3dM58QDT0pTth2pEBg
gECpnM8xQt4pc/sXVLfH8jBX8AucvW0ZgIxYzY7+mhAP5zIcHe6+MLDK8OLSHiptGBLAMLjSn7az
8fiDRPH/W1jiiWZRs7zOrh0uSQlzJq7jCRcB6AjfEAxT//jvOcxvdAS1yw7suMG6nvcv1/gU7fuR
6C+Cny7Bug3y6CS1jyQF9b0lSowA+DGlHU0fBQWllGDjkRAA+ZjXtvAuLAGQm7KhktB2A0DgXiGU
TD25cBxqx2N3JEJnL5egrcq+eWIyV6ftiyA8rsDQh6K1wMsDH22mP1t0xzFJe3oe1O3hdQTML8xX
mUoMulo5cPA8gI6jSbuax9mTpFAf33X1jXGIBAcdO+JIbWpMsTKahpU1EVJRkb32k7da15ltc9ZM
s0bPvIS3hu9lzUyOxzV4ADX8N6V3HOnIjrFz8X5E9Yn78hvLw3tzKOTphm+NQKpFU6AjkTcKSHnM
OlDcAeRSGcTBoX4JtaS3KD6xWE4v+HGIF2MCsG/tDPZLPxNeL+O9jxGG9ivMaXGrf5YuuHKUDpvR
DdBOcbrQmD3z+k4IGb9LV25J+xhgUlMeCRk5NNZRDwoybfwY6bM93gPtQPF8HS5qgr01DyZhtrEM
uA4+PapodhPcjaUkg0/VtZFmfQYDYxrKoYgBV+AmIyyF8+2dGczUp5mZiBBgChoyyZ7+jH1tfhbJ
BXZDXXi2/83a2DFfDl/AgiJTezY/1y771lVxfcpV1XW4uN5hOnmVZYmUSqpnID3V3l/5WP8Xggim
BYfdVQb+hqaz5XZ1tUeD8mpFuTGO2tIqcbkzi/MM3PLe0XG4ZRWKvUtHWVs/nPDvbOQ4ThTHB/zP
a/Vf/xGiN4jhuqorDu1YPN6+vY4GrR3wCCRdU/FyqSqinH3XZVx9cRuV95WCDGBfOeqwzaZRd1It
HGs6CRcg2iTbKXLP6QABhexd/NqKIS9BjAoBlLBNyupwfY94bYYKpZ+v/hpEB/uh/Rw2eQ3DZS1Z
D97BJfvM3gijHhJxAIC7N9gYk1m5379SQr9R7ASLWHpaXGWS4sF/Mo9uif7g9FDbGwQn/BgRK4aB
6XvbHk0cw8rLtw7nzJTo9CqOcfT9zk21QCmdcE1YxdubQQ6ZV4KRQe48ysj7Cd/6D9i3dvQik8k2
nF+H2t5/ja6Wmu2qOec5z8Nu6OwR/hgSRi9JyAjzG8qIuAvSCChlxSNKx/PYeAc5GYIKl0Ukf0Me
rMMMJ2zwOTPPNUojA0QnCZqQ6xCuTNtSdGyU7SR3Z9yrTayiJn2USCK9AG2KnILPfraXEJ6Z2Ha4
V6vfKuxbo8OrtHXziBW0EIOUo7nlbILK0JczLvcIPq0DzpsfeyEjZuQFzE8NvVcyLFycMmEqlI00
3emDUFhkFhCOuQgxyskaOxwIln2AoHV+VAYTLxRJghjDyNiLoUucxX6LC0DhobY/7wlsEbcR+s2z
XEO8XcxxkgzXTwl6FsFfBlMHZlakaDD8HbffEw+ZHDNrwK56hpfWe1naLUjg9/X4QPR9CKe2D8b+
bn83cSBcMZKus51/Ufjz/5mWCGEtacd4ZLrC3DgDjjehm9+5faVIsdWHDiPMiW01rsv0B/EEz+1e
BYDlfTaxooxAGxN2MGDcmTl0FedvycgMj4jvcRiQqZlRInxnSF7RbcQt9pRBf3weTmYFU89gxhl3
jE1Fh2ndjRiZ1ejwKRGcAq8G468tka2SUcfYOUn9TADm7d+2l9ZvXPbx6I1TlA5/CQQwx+jRAx4m
pp6Vw6A6C2+8AvVzJjDS99XjShLiJI32nF/VSBxMH2cbjailrxeQMppPGXynikJoISNBy0XMtFsd
HKq/WFXiy+0USdxDyWPsrzipQ0FmbpuXNG00Qn39twAwLc4J2kvVAx89lqPlXEkfSOT6+hPxnlQt
1WiAQ/6Zik9yxAowEzCW+x4Y1AEDhJ4wQV8t/AOHZicacWmVGbeQlkgn5s0oihaniF3E5UzWCSKb
8bNhLwixp5JmwAp5YtA5JwsDuWv+4imoSMj10LqAMKGem73y66uv/13HSldn2mAkO1qoG4d/uy/Q
NrvJHofjFg4f5cNehgKWrqg/2Mv6urPiwxGhnZlTl7t4fh1NAOFgYVPJ+IfmGLRN4+xLRDzYzc/e
2B0ftRF4GYRqq8uIAFeChdxUwLCdFKASDVgA/rTM7F5eMF4HkykBNmOIFWnkr6hUPAJNvS7DlrTS
Wry32PvfIiDQ5f9Hx+6DDf1os/7mm5dhTSTFQiqoC83U8hZkpsntTv/plOIjG0PvHOW1G6r1VrwN
xTRaAxG6HGk+ULqxeHRlRE39wUQfbnRVeFM1uwtDfpaMTqVqhJu1YZBaTBlN8dLhpcvk69IvWaWP
gVRh7USATZvXTzXxspA5KVBmys9wea+o5NPMibhMwaim37zdCZLp0jjNXwsn/j87UtYGOIWng0UG
VVvjn+1NVhLuaDG6EPY25v8oOIh8t5CkclIf+CBviXr07eOfIYGucNfLhE+Za1Pshtd/ay+HMuqu
vbxVthnqJHpe86qcuzB6LmVNOpTKFIPd15X7yomLQnO/tbqPdCjyW3dqbAtA8RNNIXxLyAdqn73v
syKi3JXhoeOUaG6Hl/e1dAJbW/zhJ86Uk9YzQ4WeE/kBqGz9sK3A7pFoydLnOj/HTjyjHkm268rC
uvu/HfljR7EyZxWFyEWE4kljuy3RlWSUWzX5LP/IWO8+/zCrxfTBwUx/UK4m6784OfGaQ7S1zb7e
yJFsL21wBMy6LQcNkwd39Mqxg9dlt+rc1+yQDIU96Hd7HDYrt6jOG62FReoiInbvMv7A8bXrWQ0k
fAKJSOoaZd0YBfD/h8hHukNIPnnemgffOw49HKwiRW3M3p8SP4y2kBMyReuMVzWvheG4qvoEUu6J
YlEL6CSPq4Bw4qFvbBF9oI9fQtAPFC0VIPcljWogu5EHOTR/XFaRQgv7L4M0F/pfQ+aphps7iPc8
8x7+tHmwamonCc/dPfjuhWX+8dCrlhBD42o/mQqCdmeITYDA01JBRIAPYH7toVntqC6Hkv00ID5l
AzKSByLPeyzn3RyfVegP1WdMeup4XWE03Tqjwg8GGIPpx43lXLqukrrl7wdj4Reihdw01BUH9YoR
M4zidond5ZAPt/Pt1V7SsvaZq+E/d+cv4+devebgx4cSmiKhVpByMgWjBquLivTaIRPkpcQmhMKm
77m/D5Txjy6cnfbIHQup0txlQDuUIFcXxsKsHRASUFI68LaYWWbz/SHf1RfLJB1o0zrcMXZAyGfX
eJaNwJIzekoIh9UzI0cXpj09PyRFPVHqojMffM+WxlRKlXUlPWAUnYFqJ9y0AL164ary6wBwfAbz
eQb573oJbXzcdopwYAxS2Ppr7hZAuOUe7WZD8d6vWTEsW/tNzKBXxYG7waYOz7i1syRbdQmrLWll
oWwNZUKhpoSIdFrfvMRIwUJdN3ZNNJzevA/RGSaIqs9fPbt9FocAGPi6CVktUu69RyEMsGKO6kvx
wzHioWC1e6RxANEDDjEl4gF8fm0f+cNN+7OMz1JpNXv7nF7fyphEm38J+r2QDJy1IIZlzOtsQeS7
oHpHXRAkO2GIB4plMQzEYapry6NHA305sqHrGEilQ79vC/b0RYIPsvf2YbISIcswQgtMYCTTSLbb
DijnhyfwVnPRlr/IO/UuMRLMnDXIeff/SXPnv63Pkpt5dgCbUwfpeHN/5U9DXYfCq7uhLuGZatHq
N5KOVnRgHhfBMFOfrZUTow5mXLYKsYWte2xKiDT1u+ZXBHjCrA0cRFbwWVPKDUvTprl/Jp77EHbR
LuwkntVkkoAEcxXYZJ7zX36b5fItlCtBQXi40qD3eVCxRRuDw455H9Qfb9Fu3Dm/6BuDOlLg7Pok
B9UW2Trc3uIfKGGARVVgS0+WAXLhy5408tCWkjEZh/pk/coYI2YVd1VgEvjCoEKV5TlwBtu48L4j
HX7HIeITTGLpAtYuoPUJpvr21uHkjJSoWeAeRwk8ZNeUo0vReFqV/7x9WEyYH53hrsToTeknjg9y
osT+onwkpnC73HciUSRwPAnhB2gc46NXKOLFjRqwzlpMcJd5t3PAnpW2ULdkYeMIjL5iC6Y0l+y3
dOMjenQwfFNm74pREJJe+weAYxmkhQOEf1ao89PZWy1uxyVZg6wYXeJZuGkHjWwIFZOrwhu6ncJo
yHYakd8OApfjDKiZ5DbDYup9MNHE6P0+6PMz9OKXXlIxhqzgreOqrhc1pBZkAZ27SrgFy+SBOwF3
I3fV27JcUHqslzEgTr3+dk11j9wtODmeZ3dgRIpHaAxYZ8dmafd5zGl69qzkkkuQdOasYPrNPuet
Ep0nzxgU0Txz/FR9XlhUslePR31EyzneVKeHT9+qi2ZCifRF7H8OAPZTuPLFVo53RDQFKM4YB5vI
6KhVl3KvXLDnkx+TNAN4H6R4lTURnIJDRx1q3t7LgO/v0LryTe1RNh6fEnIULQHfNPC+QHZGLSse
LTEpY0M5gPSVkE25IO+ysy7AAclCkvdSF0sJF/QN3dTFNMSduwHyKFXeJRyqnmIEBuT++BANcjSH
kJohcOkGtmg9NQ5teSgudTgz53bOFa89thkS9cWbjwStsN5eALYL9iqdPzRNwwvOEnjWDlQdAKOA
i8sMzgG+I4kEBqt4pvlj1lGYTOl3Ol+SGagNSKJiBvW34ZRUT4nEYUoZ5O5ibZY0JkE+z2pwdj6Z
4CrlU6qa1bL67iUcG2vlecXAHq2RZ9Vw+zMN2L18AE6rZKcaLFL4aJ9tf1XU6Y0AF0WvtyNsK72x
2VLLMrulMA0CAlpRPaZ/BWfLaDEp4tQePkM+ndMIlHV1sfQ2NiTNk+i6eByJh7O01mdw25Hbyv+y
ZppJd++bombE0lYA3mTet5R9RQ67z5wrdLqjy5jfnfZSRKoXeKGySB9lheEc6jhbMYxetQ+wjrLE
PHVbLIh1Vqzbi2rBFc8DON+mJdGwA+kl6aBJCC19eyKxI2VF2kgIE/loGR4NhfD880vHrxH/SPdC
JweoCi5c77+7KvPK4hHcF7ein0xgFzVxOyUdwfm2pLQGvOCW5RWUKajet3slxktMNwCPGy7PJN2u
2donsCvTzLgcjtORFjXVmK3Nac9MHgmEZ/H0c7xVbUgwIPQ0ZeG8b+4ypQzbORGw4N2Lu3wL/LDK
uy50eL3byyQezZdN24cuHgpVqA30vfjHkRZc3vCehg/uudIdov0W1xO0ERX5kiVsC7Wh9wAjIN39
kyX4+09y0j1vx1aJpk8hYHUSvZXF2OOasyiXyTkZuO104IZ2unOmHc2FOwK3mbaWzvTG11Q/4Jv3
8RX+5LscCNBESkQCblx+iGX0frtPDt6G21wWqthtSBrYkIyzuRx66duScvfaAl7SXXOTH3Uv9+J3
/eY2EwSVouxfHcWRM3tXiLRQiT/t0PUlha5DxFthC7uIvpXgBwvpOiNhDjjyjwllmxRGmgbXU2FT
pgo6fgJpOiahqzuhanw2SMpb3Qa2n3QrxudxuhMr1b7bk1L2BWe5F3cbJjnkEb+JI53poVufMYZC
NBw5E+9KKtL4zMnjKNir/idoO5mgLKh3FZXl4387sW4f3e7E4/sOXzWFIaNQJ0nKnVhKnLdr8VTA
kwdIkocVmr9oKigS2EzRJYaO94ihStos1vwaxYxXR/LPQw7c8bf5b027e87Fu3nOU6/eMmsdisMJ
1+HvM4eGTGEuMRrjfvZCPvCP9ZpMG75i4Vvi6qaB7TfWlgvHyXOpuyO3UvBK/ZZ+QtsuZWACDW3I
JIiKouk4qo1CYzfw/BuSisBZxeX0zRG3SeiVH+F+7nKpJJYDN0yGYXLNJebetlMgVY/tdnDrASiM
cGa3CY8jz6Luq9VjgYJnitqL2Z1fUFvcDcIcAeq3amL8qcuJiye+Vz+zf/FMjM+KLIWKss1KiJFq
99hMdg0Sxr/S7UBY6X+0I/+IkCvYCZXC6xMKvTiI31mM737UV55QNVsRrBFSL7E5LXcg0aMfJQ85
FVbrn4pFjt80xD6VrELByHcmaIRCXnXLn30xOaUjwvyJmv0wrdzE6NY1BLTrmVJ4hhdQ/Z3j2h42
Mxsm92DCKEgIe6cAXxivZLNaPmSzUP+W+ZlguGnz+lFsqkU7pUAmvJ69TP5bRyxw9YfUKxLL6eWA
a4JqvjRIA8c5hVC0NtUioCl256pQpOThXvSitq4VL32ENDxhp2rLotcHrhVpr5HHTEV/nSUJZfqF
2C6QewYjdeNdUIl6Ov89IkJJk53CBFeV8XaYzj2rRf7FaUk/rK5rY/Un1W4R6ITiT0Laq10KvvlZ
9eH2gtFP7FEWwHNZ8rxi3Sns6SEYLJCOgSmSwiT0Uf+FMkTEtcJLMN7qaKiaW1tJ9uOgsq4mtLfX
cfYSrjxTPsgl5vOumG0mRsMLiDJDiu4YjkuPATEITtMEodB7uRYdjODS0QNC5s+xiYSJKp+TEhTR
weTZ/zab0RNtXbk22Hai4HoM9zLEb4uLbaFsgQfqPpTgK5qYIWjTJnDnVDQtHZkmTEmmD7PQoimg
WL3gJJbV/dBBP49t8DzfY5bN7pLCbytorN0EhiUgt2m1tMhy8Xim503MJEW38I0gGsI+UxO/pjMz
20hq+U2XeiL9OpcHpVIZzbuP3Vpr25K56yACLNMrafLEYE0zDDE6VyCF8u1jAqdqwYmW4uUEA+T2
mgsazSnT+hRQXztm/uOj994hhR3EvmDYljgwIW3tGvxOb1+JyqERwSKx7P5Uu7BbLkAI+OSMmmR6
asIa4e403ZzYRoWyLz9dTsnD+0V6Bx8oOpgSRG5F3l8h/c4zil+1HaIId8CmRuPLGUXxt0nxmmop
sh703sYMDWHP8s0PjLCcpeFRBkxXO0qJ7J9MULiC+HPWSvidrnKhmAK/r4YRzFOmPRciVvsS7fF+
RBqdnhZnO3W81MmUGyBduBg9nHnVfoV9uh9dLUxabIu4HcN34daTNOckYyB2opK89BWJ2KI853Ap
oo9PMF/3XKOuiH+D8SHR2mAcTChKsVk2OCWkrlTm/bCQlodLmaxeD/xJnoNl4VXXQ0H7sVHlPpz8
npayFa5e6Z+q6c1nbqYvz8OMjiMRJ/lzhMBukEfhTXZYJatEn+97z52cn5LU90ES1iAqbfRfwSp5
+YHvTd4/uvLkbfl1/YC+u+TilGauJuVi5LJ/uWpMd9ZFOQT3CvfW7i4FzCcfp7ZX2KoP46JuHIPr
jW7Ya1hmxyyJRvBXNqMB+wjcrhWpVi3JqygaUnF60pPRsL/Zb2V+tWI9hPkEmU+SbAAc7Oj0omRD
f5vhu+28NJ25izxlbLopm8rTFeiOIrqhD3Ivn+XcXaqNF+ciBlxiZ/24ZpafVSBM+BLahcCUwBCY
+74V1BpGy9MIZWcRPExp3Y/tnECIokC2lCIJMNaJBN+fR6gk2jGNVUXLRvXCv/tbqcTrltrUuA5W
3L1YNSi2hlkDYfOll604FQ83rseCFhCSO8spUejiwmfDS9z8ktn3W0SJA8SBynCJaLnoXET/lhpY
fiD1OJyb3VaNTiPj3N2H/490U7uovuMgiS4QEvcuQYVozmRJ1fgtET+0W3sVt1thKhg7gDfIRdxm
iyDH8EKSEAW6JcqEDA2Ng7vjLifjjGdAQR3Tp12QoZPjxP5IdwZPYG7x8/1vkOTXTX6VwYhCGMgs
bg6c3xU4uQcuXgsfg9I5lzODkfeUcu/7pBkJuZBKYSmUUUADh6y+K7faLQ9xoWbUjsvyFUHZcCmG
J5nu3MTQ6bt1SPFXUsgzGJ9wKbrB54osET1/QhzvbhGPzMSKoHCPRAvo6/YtJqaRf5J3leUXwhMb
vpeYks7ibiFQYC9qAaDJ3JEJqtF0W4JoWCaG9QFw5hr094yfti0CAi/L1EV0LnVb6ox/x+3PBdS0
GsKwaSUr5AlwsZpwkTnmLgk/R/QX4KtYt1DxK6KmLu/0GjAkW8bCMQZB2ytioUJMHIDT5dTL3Gr9
qdGjXROnvN+gRvS18ERlPzTsu7GVNTDx98lUq0nyUGdpdW5rE/g904TDMyEadl5Qbsfs9STNbu3U
cWm71eU272niSdnc36/1bB1P0HXVGab7VLpyrlpLb4FGWvytA77MGpBRv+th+ZDXr+Gb1722tcqJ
JYW19d9/M8WMnaB2DSQYjaYdy8XJ6EkRJXWqpj6fSmU9abT5ZyeDmgUCm7s8jn0Viy8MS9nJ5c0N
v3UC9DjoDPXXflG9eU2ZmFrHQId18imi/0vUhgVdGyEDlpDLOk2FX8HH84Y5i4Z+f4I4iBVYUyDB
JQh1D3JG1RpG1CMD/VI/SGAwf418VCuKsAH19jH6UZmQgb32XW/m/vBpP5T4T7VwndscHdNY1Ewr
FifJaBFuJJjWEINpKTADl+z4a0A80aC5JgQHvu1PWFqq9WTP0pRmAsj7Lh3mF+Ad5mgZJoJZLING
Oi6S7yppXabuqSAAbbAL/KvM2OiTQ5ur7iE8H0szGLgTznvFl9zVxcHlgaUosTCT567GV78H8bxy
N6ISESy1fnj1ZoQIzD93+mD31bF7Ucw6cENeruAmwrEASdreD9Lk4vTN3sYJfnQv9Yrj5UqBTWod
EUCa0WRKN5t7rY26hINA1097f5aNbbdA/pte5tPHtFcKGeVs+whE2PyGPN5UptmjMOkSz8Qbs1wo
GqDm7GxevL0XrHMTRPsw+YAt+MwO/spGKzjuRoQr4ZVFni/67j2n+gvIsVOd5e5euuHQx1sIv7Dy
0hg8Y+GWn826QtMb7FURCjGL2/xw6PyW1w8AGNqYnfJ8h1LqOYKcjpxwIWaCJrRuX+70336lH12Z
sYyQno+7pEsl/2I/0gfMhAYGc9Q2JmLUfDhX+1WwkKlnrgkhLTvY7m/onCu0KhHenUSKtbB+QaEQ
HVxwaJ6+kPlHxXA36I1T65t2qoZ/VaibRyHAnRRKEKhvZsNpD43QE9rDCPuK/FB6NXCDMxNNbDpr
jIuOfgIzRIEInS3w8Vl1AazvxGahRxnUb76zcf2dWL2XWE5fDHGvwOLPZVFsFlG/vVBAsXJWQvZD
n3QWaYKqO0Q7PKZLaVp0fBMwhW8k3fpuaHY2oXQrQCHxF6U/b/D6NjsEgkoR+h/WYXsHNBkzfCwM
LnqoNRBDvEuXtPfJVB9/k3Q9wr3Xhl8ZBbnG0a/u+HZpB2XUTuUmwGI81P3/IKa9GNG6lg+PTaTo
o3wICbzJBEf7dS2yKQvb6lwnhNfwF1t8a8HeA5DN7Q/81TKGo5x6zY7/MkMZqx2WRfpwVijq0IMp
TMMLemZya7htNDPpGu4Ut7YOWVK29T6OL6gD7W+02Sq1iSgRM+tLy3V9QsgTVKA3e4Hs0mpqcdSe
LljgOX+r4th9eY2zUNID8vOajl03kZwxHHTxxAsg/LJKgBNOdicNYxY8PRsjSaOOPh1vZOVS905B
iXXygGyLlK5BVSsojfP4AbRog/3h1uTsYAPSkIf+z+3Fm0abtlqEW9A6q/8YtrP43x1GTE6HCoWI
fsCS/kgdLpY37yDkyfJU5a1IwUKGQOIuF2/J0JGmExhMSzx4km6fYDANdJj9sBhC6lic3vyYpKra
6RVa54R42D96T4M8Pu67b/Q30mHVl+M5usIWRo1RiXJp/4oJamRLq990YCikOE99/ABR7o2k8/hj
m/R7sxAljhFZzeSUkcQmEh7AMwTrEVLIkTvfIuYO9yrzZFTlrL5b9/ZAdSMMPFwiMk0M12yKoWfc
4W0mSxY0nJ9K4qc+bPWfpjbjJEy2wOkFN7LKT6Ok83C4BSnRsQ0NPzeQy+lfMW9g20f9AY+jJAYN
K+mmEXA8aIjKdwFRpUBGXHfcQ9iPUGdfCHM0RZuVf6YUV2/qFrClgN7PQNEVCo1y6QiaG71SbMIV
tyuxjfwxP/AHl3nANKRBTwUA+0bDli+4amRVcwOx7RAOIJa6V1FX7NDNXowSbqaqhmz+KVGNBzSE
seuyaExRS2EBcgyYg48V9bN3wgBDHb85nnkwOac4AlNkh7bnNnbS4EU8de0Y1ywjRNq87NeC0vRf
RQyhLhqFQKmgywCdeSPDv/8YC00fK5t2B039PToVdYyZcr07zFkQo8ZPlO3dqFt5DoijDFf0uQQa
0DCwlmprmW0u8AjiO/VP3liGL1iE1OCsA9eYLjZzrwOYcXB+b/pkx7GYjXMp4qqyEHW6jfPU0c0q
StNmwXTlaUlCYq0Xpq3ouyrD38iMiYzNUy+u8ye54WGUG3BZkJoBBt1hpzmLL+Y9L5TqsYMqFIrx
9ETci/th7aFOcAWGUh3DYvLftViz3JkLX4DU1WONCWnEDSK7lxNb7PJXE3SX+0zNB5EwZFpuKRwN
Ll3/0FFhSHWQjkw4p3OPhcjH0EL5s9s6ovN5W+HuxDGj7iCepAvqJUm47lWxnWIJy9bj/OkGqgXA
NFwJJcinuY41iqerUqlZQYOg89qVAtbV89LGPmw/aNxudpJ6Nqmswld0wX+fWHyVokmdKr1r3Yz+
ZuMKkgISYvDCRFqdiAVrgp3ERSQ48Vf5w9fUv2Hj3TjSR3ijNoyFqBOqI4vZzVCQdaVaD8KX0zoc
o4SbalCDRegM3rk83En1avt4NFlZOIoq3BmcmTKzWHZ51Dwn20QBPEFOLqYLd6SkmzAXmY6MISHD
qZZXIeOAwldYK78htiSo13KqBy4CPh/DJZEeMWkJHzQb8TriFY3CY5i7zdxsMrm1meqxq/P8b22a
GaGMhqqL2wI9UustZnIHYGLxD0F1/ujriYqghk4Xsg/k/tG/4D9PpD5v/WNSIiFdgr8eJ5iOhdJy
v1GPHAcE0FE8yyoY1T0q6DD3Ngu06Lbgzwj8A6ra2Iokh3LdRxN9WyO8AInl3Hh1Xj0z8gnuZjKI
kLFFGSbJMeHjXQC36iJjpfx0VzSK+wu4hbwhez6REtYtodYNrhqWucL5+Dd0wg6ARIFWppHmOqSO
Tgl5GE9Lv79ocoJEyZfUvlIIl8Dgus5QF0opFgc04ZJ1Mq6csMuySfrXR6I82Kgs1rkTuQ7HCA4Q
3Kw6wVaRb66cuEvOtQdQoyl9PhFN6XIuf8m7jr0XZl2WS75/8Uoe9pvC1905TnyyhiwbwQ6QtSn6
2HMcis+v/CqXmeOvNIOx8P+icHEbIzoNCnvUf0uQZ1uCyfP5QpUy2nm+T2yKycPCSu6IRUwawb1X
VmKX8vFQ6r4hLJ/hu5Y/yZMLFiI4kcbg5PLqb378flJZOF0520tzYobsac1yFoN1Xykr14MNdCMt
IjoCjlwxcen1SmvdO8Q+FYx8fdjKCbPdNx9KB+tHGtZqC+AYPmSHNeeGA7AKstCwpd10Sj0WKOZC
X8ufU1lbdvdAU6gFLxqNNJqQPfuU3qe0pHSAyStVjYEAuVPo73lBjrL4rjxKeUKBNOa3SKqHo7Ix
21xy55jsF+suE9CIF6jNgjbg5IRwJDZ8BDxKOmvM2SM9jUG+ez3AzGuETvV6qAs9X4B+rBu/bLrw
pMSBcWI/a+5Z4VIj+/EzCN07veXty1ySNSYQsj72rujANcZBdKSpD6HglS2M4Agb1oqzBmTd1PZO
jqi4zTdtIGfplFZwo+0cg0v/Pn8OEAwakoCr7/BQ4F1OfIsAsSOxxZPcFzVsTm8xxbpKV9EqADKn
gx73UEN2dFvW0HsZ9GPMxQ148NTvW/UyIfFfHviqZK+CIyN2Wv6RUFVsMECR6sm/CClLfUiaOf0J
t6NhPQEIA6MPkkpfCxrDMNkjaCRyQ1ZakG28XZGyXMPf/9vR8SldbtHIBbsXNSD3NZlovYPzQ5QW
ldNkLXJVSCDqYV/GmLNePFACpCTYSPzyfFLIE3p9JAyL4fkTkN0PGBuC8A6Dt/geG/Tmmisff7BB
GjBNOXwkyVw0kDssIzaEKYTYJqLo5kXhhLBqhVX0lilijfwmFLnMy59JvLlDvnDPKBFAhl+MyY4/
alKLsQXTfoB5695ovxDgbiuEqOzzaA2/Z92LAjbjBnCnrk2NMVE//OowRLNsBgM6unXdbLuUeybK
1bpjeJislMYxfwjoBq1FcOs4/fwOmRu4bxbv05KkogrXsHTW28wp60GAnUpK3O+CKK2Rf5LsWvPJ
S6vcHAJy9PlVahGMVnCffqO47cilM5O5FC7qhFtiGgwhj8I0487haooFXxnsKRkln6uqmfMyht0U
Hab9W+jxDJumhLeADOnnVToKiqXX59s7/1bw2lCCKSafYqF8YtznDB7wNeaq5v0flQYhCAUy4CTJ
zbiLThzri72VcHn8lpfkdd1pRvjSDxsxujNv2nOrcriUx78gu3R1aPjg0S9aZo1hfEe8WoshPwhM
9/tyegoS/DBXHLsBa1gYFlCkVn1FayviHC6whxr0A5y66HUS6SfPIg6njr8X70CXnreYuWBXaAMi
XjT0F2I8Pw/y9jDgT4HxVnnYjpZmtC6nKg4qfbFoQlXwwnnB9knwMqU6HQIdR7ZSvWPFuZXDjn96
wnV6JR/SihxTN5qQcdWSqOjentkS/6W6JZNRq9Rbfsl6nrK+zJv60y6m6KjoG9ucDDIaWBp/f5rv
ZeHre3zcaiTDYP0tSp9XFf3GvEpn5UjWIUq+iBeKhCQBaMJqpX1ClU3YyKTVsubx5ybZZVPJzyCP
G7kIJ6v5twx7nE5pFUeSRC4le8Cw5cFpxeDWEzMazU+qkKWlZm9GnwAXv87jlkJbsPNmlNzlmZQl
lAgEJK9evYOmxn1cWQO53MLKhHYZzVWdas7kVveqD8QgSyhLfqsczNggk5iNuMozzXqjnasLyPbY
82WM+MaCn/gB+BWxCc8RDi0VayHrnPaQxSgwB+XvQzMMx6FaSVTYKRZGG94AzcrWweXNEUL8qyQP
9K5GFHJytyr0cghqjjC4cxx2M8vmQzob0uWHucPTqLPQyFQ14N9uYGYjCp6raZigWz/pRqOiNyr3
Wa5MIq5wXt0M+PmFh8bB/NSjqgu3eIWG2RWbCTEkf3LlbhusbDYN6T4KyPvig5Q0qXDs3NjtOn6d
3GtkQycbDGpS7UDnRMW9No5dDFWmr22jQqxneCQPBq2SWH49NH8u5r5ZULVFBtc5QFGMgMfF6AEj
vAM9BAZbsqk6n+5AL2Hnj8Py3LSzGTyQJTj5AGjmxrscAi7KS7ICSTCLvqk14h/T2EFXYr2Q+j10
hh0BbLweRKLuN4TAeuXk20cgsDmNY9akDEjRdNK4IFAXh/6oxbQ+NVXdsRkmTkyJLCeX9a5pAfIC
Q0u12jXQ5QqEZCcP709WuuLxoX3sn1CBhDIGP6h3P3Qqy0ohkabL6RwR3JRb+Q6OWgMJvtsk+Fpp
CbGfOdonUDNpMQJqOXNXh4gO8vKyRqEo7iH+0/wxy9LM7AVFynN3QRPlu/B2fUqfgmUcQ+5c6/Jl
GlGc9CApX459qRxYW4qWrOQF8XydpURYd6zMyY1fU8ebW841fPNh/GwL2/aSpdnZPnISxAFN78Oj
eNOHkBKVTFIX4Cl2KfBVnfR876Jwt6MK/ZHeeVmAUjVpfrvOj8F48jwo4MV58Ib40xkt6YCn1mL6
stw+3WNjbOwV4ilqBbQ789zG6AnmNy5ayjuK+bxKb/BSpXJEBbkqXyBIi1wwVqfDIgN4Kfzg/Jrs
j26oQ1Ft+r+7eX04Wda6l9NjMjcGQOD/Z8OPmuS1aIA5sbkodmjyRIgrHQ0kJsAwOka6AZxSvv90
t4OkNbDveHSjZ3bRwK5OauLWRhzruXN7JleXuuI4ho6cAFlXJO8vsM5V4JWSoTjp5Ivuvaq/e8zM
si8V83RooTuPPwybMc+KCEpUjnf4Ft6lKVTUPbRyKOCFFXd4c6PbMwJbZ8yy2Q/6FCL0M90tFMro
ZuvY9omBf5fBABiEPVNZoXRyTz/RsKh3Hp36C+SuAhxJwVAj4pxTL040lsbGX/awc2v7breO6BSG
II8ddbXPf3v7OYVlD4IgkOlyIAPOAbP7nr/HndLrthAeLHbNH7SOW8mmKwBH6F5uMeokwRXJCmNj
x926bnvQ/dEAZmRXlMya5rQozU9buPWc9swJB2yfflsmY21wp5/ovfHBSeqe0hlB7Am1275sq4Ln
FPYX7uerMRGFZBr7d+XbASKf46jqNLJEpRHBuU2sZ1OS2GIXW9Onz2YX+odn1/qwEMInSeUD5bgP
gHH1COxt/AEZVXDMxrZHBjl5uaFpYYIkEzbe7xO2sxFQNb7+tdK8NMFf7P+wnpS4GXcowpcSYPRI
EOB3IL9X4WveSySTmsSOrBNhCprImnLQulLiJyqQ2/4W6Cs70FTTwDXhvC49ZerRzdcLcQGI1sxY
IYuwjx/qOybrDKWTuHzCDXMnd//ls6NKxf2D8F76dvFbI2Z1fq7oCwg6SdWWsrv4pLOYUQo5h0WQ
lkrQfWie4EDLzrdo6N8A4siygTGeedO+sdTdMQUYHecGKAR9fNVnMY7lOGE9/2maTUTVJt+qgLYO
6QFl6MPrGrTmYTGEiPdkk9cXYPVUWtKhMQYYqIE6/vXuqQCY34djka/g9CCJbG5HQAbqcp+eXEjw
v2MbdWMKxcSpczvTKMsZM3IwCKgsXlanN5tAe4NOTr2NEysiervSaCun74mEjcwijE+DI3EjIkEs
nifUzBz9HolHfUjPgG/L5Zr60IeKBj3dTaw/9HtArrYl8auKblzyIfniI+iDnpsDtR3UdpfepFPj
b9FjPbfqVoV8Nw2RvFOSH/x2OIhFP4fc3kmLmmpPJpSZh27HC2oPcq4i0NzNobX5lI9o4JpyKKxr
11zZ5GB5CRrCJMe0WzPVm5mtfiFICLHamsF69RDX78GUaMiVkkX1lD4VJG0GDUnJQcT1AZklDfjf
U5Dnb6l/tchtVDJWp2NJZaNnTKPTJIOUhgXF0hVyDu3VtgqNGi484Kz+tPd8gEbY030GDgnvPM4L
BItZI2X/haPg89W8jFS614+T1NCyl36e9oSwEUUvfjKyd/13d3DrxrODHHkszmXNWfXE1rceiy4r
YkIQvl/+io1044flS6P/ZXytUoBZflbw/0Kmhb6JECjwe9TtUg/pQzr1l+IqOA+3MsAmj9f1TWf4
/i2L2/FSk8Ns6m8NZRrj6CgHx/Hq2/f1E4mmGoWVIM740otRJDKOejN6/a+kyA5qOD47x7Z74hG8
vF/0rhf8C/UP3Kz1GyxuYTvUgPO0IUWObAwqWSUcqc/ldePOd3Bh8Bi9lch7kTXVWa2kv+S6Mw/n
hb9hq2UvAgYVa4dPImD7MxoIGBetMcf9z5h3xuxEe4csKZytCQ2mI8KE/wmfbkXiIaR/Zu9EA7Vb
+B4OCaBiUn+DM7LoaQaHO1lHdJHfUhD/cp4gQhuO4mEC/TcDlQM2zzgjS+zXSyBxfiFpCSwX1+dG
CACMAClAsZly9haccLjl2FN8V5h/nr6XbNO2/n3tAD/SO0dSeVo4pDhl6B+1KbhY6LNWRYWbcd2u
y+Z8qWYxKLo/SlWmpz4NIJReM3RL4PgtYkLNEDtv6w1DSp/c4Yol1Osr4MsXmEwBKq7Dt63dbZaq
xipUtS3gCuyCy7m6cJPUilO95U3IFC9o8ZoHZTZ1qJC1mgPjfsrTPmehtvrdl1ObgD77El1SU8Wx
ZNHC/4eIUt+wxl6mEX5YDPjOC6jGthngt3/tkm/y2hviEBdA7aKv2GQY4sEGUwWmRbdCacipXTXB
gkRnJseFgDnaxAj/P1an82CH1cIHqCSNgC9w1MRNAjyioXW2lGgxJaT3JyMI9fSjBuSZj1sfWioc
YPhKR98MqN2F+2ExQjijrE0ugWZvB/SS0cqUNi5dcGkdATmdOJgP6cyxv/NWXRlmrKpowjKL/TWw
fZcNJms72pxI6/71GOdmVuwkxshiQOivfdtGGl+9EosbMnzmQcBe0oKON/09vke1aTcXfaAaMJkv
lZx49KO/3bSFBg4o1DH8nkt39+/9A1iXn6aUfqDL4SVHnjZXqGZJoAd4YmtnTCZVAs/Ux2bbSMVi
A3Uw8WikaH9HzR62LzIYwiKdtq+ZVz8XMqiO6MpSHxEbqGNWhPXAyBF0O164Ou5GeZT9hy+cEcOl
t+Q+6XmVsuApQZMCERuGmvSzOSGZ2ywN7xHEh0S6cWUpiKAsljdfl4YvnoJZMer9KHda20ZEaPHx
fpon5ea9vfHXj9ug+vMLYrgrsyLO0cgismHg2vIFvlK9/5gFYwD/MRpc1Kl+Qd/Nu7w856sEZJSK
7+IXpJ9g662aGXfIAy5oUHnwVCh/qlSvceDjf4l2YinXLHtC9jBJmth+BNUYjOoslmbuvdKw6DRp
HnChzlB1AnmuZT0F6rwRnio/yUbqfEXRwaofMek0FQL75PcMWf6mRM/GQKYJft7tfCh2lWlZQIGG
Rez5CxCFOBORpMssYuoFnW0cbBJLPZ3KQf/wIpMeS/gRVmz25bCw4aIhCdvUA+HzGUnG/KRD6MVl
00pNS7/0QJdxLk/rvnecwxlablRuQJhPZyRNhLPeUSACQvrQX8nJRtBwBKVEhlH3SGPcnFFoSYYG
vLTAnUW++kg8TZKhT5Anp1wbyHeXrHXQbWj8mcRythfpVHYn/2FRwRHp059Gpn82ENJ67ZHuEcrh
lKevxhesZmMnqwY8MtmYMgAnyt1CF7pU9huJgz7wN/oewPFk76Sz+1zgsztLKS+ejfnzM8Y4nBs9
dx5und4LihcV+nJlq9DF0Qh/o3F0bM09EsdPumSkNnogd6bNo1hyHhV2U/y9fYck59D+ZEbNzHCs
gfSdcZ8dMX+pEycoEGaYs0mlzRIfu46AFQzZ+q6PWB38CUy6RSTkIIc76uJ3mHoTMS5K0khwt+4v
1FeZcerDMY06r8REjPi323L42N5FSxuebx4JsweXPWMmgqIWQ8WtUxoSy8GxhY0Mduu6JsudFHL6
bCG8IwIZQ4ZDxLxe8x3VGTMXs4JxRW0eIC1LzNbhuTnRsPVJpg+kp6uzNCBb0JyVBhQQElMH5NUX
34If+79eTghBKr8764G3rJi6l81YRbTa7aWZ/s0OsZ8nOqPaARoQwCRDWoBolo+BCKgK2uTd2RuL
ujz9dukrLaRe+8i5MdcNYCZLvSIFFGlh1GtPOKif+wVZ1uiY8p0LmazqOnm7AU9Va6RMfC83Nn/e
UpqosPkVCN8pf7NgV6HUZTMkDTv0mdyk5R2AD6JmdvXenLbL7Bkg1DQo02LoDzhxX0R55regx4Jh
QWN/3QB12YSGU9K8h+L75W4IC4kdm8WLL2tjAjmXS4H9MeVRrkRe7kc4Rcgao0czdnoztC6MfTMl
Hbz3/rg9rErXPFiZZSo7zVa3rr4caSLojodukzwqIMRXAG06b7PwAhNMV9M5l/BbiiUmb+NVaFu3
Jycpuc0X8WS/9JUmR4IfPYZnBkhdgGoR7DvqAQptCKiVA3HG/9oYOG0UwpJhKPNG/q73q8pTMJYm
7H71bCRggSwcNlyBo+ZjKQlLPJyOZMHhxz/4Wg7s4dDVIPgAJ07isxEgnFuUJKB6knn6/Hdy0sj3
7ZsrpgI2QkmUW0rBc5v5M/4Wc2Vj2IAD06YhztlDLv0bVbgXKlLkoYu7+YjHuWI82+5EDHF67RpU
UtN6cXU6gxx8rC7TjitAhCGysStrCL2rYVW2dq9II9TAQ0hZq51YonL3P5/YnqoeidpcTCqrspoe
/ra6KAotu8+BeJYgZz1kXd2dryYQwrC1WkjsejsYSdDpfMrCoz6QXFDb/uvi+pbtsyggYoMWM1qG
6To7uRTVPBUZdUm7fdz4CfIFWLCgOE6OOcSuA7davbOI3em4C1mtJ6Zj6b5FgBozCtQzH0fopzax
gb0DaBpqgwqGmTXyFr4vfxFLSLKgOTtCS5VCnAKLRVZ0S52yXyMvYMXu7MOZiemAFMpAbV7qpO/9
4wnSw5GY8d9nqYE5GaOEDKpR9bi+zPYzerxFV2uo6r2JwT78klEyFfW7Hcbmw2jJUW2nc7nF/irD
b2zeuA7Xr9v5aWa0hTSiIXMCGFXIJ1fTBMI5iUN79qjRebTJOKGgka+S43AFFtL7zB2kPP7WEDRg
6xkGpMFTrYYfXtx71wDTYXUq2XbJTmqbG6SpZrOIOcvGW/hFzueWWTjB3FqfcGBmFYtLY4nBG6H1
yalwPCMG7Ppx1db70/WJHPZoRvzBHBo8hoYM0TrpA0UkHcTksKwfsLTPj26NtpcQgQUGGjgnNo20
11FE4VkoQd1u8vM752Rh+ibPKnwL3ik+be3wu4x+k6bP3jslCn4pgFet/jprWP8PZTGrKjr5cXWl
Cfq107MdUneP8qAuNHMKOGmt31qr4pVBYmofDFeqL1zP4/M5h9PvYn5WLig472Eh9os4JsFMCM/D
0xDSXQIHVOuV77sG6VHHIvNrLu77EqZs++fX6gU8l4E3vnEKxxmuJU+MwcPeUWkvbBCfjy57/l0V
CHrXawDcoELzzTVhmectM+uKVixWdJIzRb2D9RQ9zk/xoykpFAbVROrh6KaIlgrxgQY59oRoSZ5+
YaiqJZoGKJFy4oB6KEEAkVDLJ+EVQ5dtwRFue7371fye5LOIW1io84GIqos0WTyFd3TzlKOR88rS
QQxiATnm/pvugbCI91lpw704Cd5N3wsLXGgq7dMZojF05sf8vLCIxKmgox8G+Xi6HUzY6A4Vr77F
keDr+7Wab3716d5OrXRPzJxI3MyUbWONKdnnHVn72XZCGW1Tttzq7gpA0y6OrcZGC/1Kw1A8/zQ6
XV4IepmIr6oN1sfFKVqbSLPyj/LhNmofVjYz8w9z3wYi4nc2k69X0gdfu5r0iXvsJC5WwXSIPYu1
UI56Mzy+PFSernijah5Y4dhGQqSmlX28AkfchgtD/kOosblYQJNPWWNEz36LaxjTG1uf5jGYsqEA
t5+aLyKr44MZ9tA0y52hmKzdFHL2bO3nv6u+i50a71sSa7uMCb/9231wCzumqea2OYa7TUHH08by
O02Zs3jbHX/AmWYfQjusl44uzOB4KNxxvX8Jqw8gQQWrBekxsIcgSrtbpp+zwfc653A+mI+CzNOk
4KqLwKVrpohBnRC9ez0HM1jxiYfUemLmnfAH0Ypp6s2jSXkRqR5ioZBJro1r1sm08325abf4fDS9
Glhjg8yCGc89D1oxXztmGP7Ta8nFJtHa1j8szeXqdS1cwp7uVg/jrIr28gGO3lsu9JH0uPg2QsCm
B/cR0Ur8HcMSW+8MSTfr3g2yiuvxiKyYA4W4sp1I7xi9ZpTTiXG8Gm5c09kNtjDHtybbgVhdKL86
5lSG8PKcFC6O7wV8GuHyfxBtUIMku39ri07wk09yz4SI5LcESratTCb2CtR5h8ja+tJtmzJPL/Po
De/IEF9DwEG6jBp7kethfil0qfx/U6dbouNCsz0wqqNkJjYVMPrV2SQFCHtKXZBrFLqz4ksr1NYt
sh8b2a5dVnmLh836SjCKV0V8BaiURQ7KJIv/SWhxiSQx/iJ00QedI9iWQrqdPTypOoMuafjHDrK7
4QLWLVErgB6/Iraw4OKpkqcd1kjmEcgFqI46P7HkwDeYyyBeUZUCqiDsbAnotyBEcaiZtgwflXOF
pp4T4dIjtY2t+ROQ36PP+GT+tOFfpI7jQ+IqFKfTZ5Gwq8sari4aCt/dP9awA/xSMevHCNEcbHIZ
SvetMxmJMtM+X1JQBMhPsreJISxoWtt2P5tYFgb98TpzruwTd6LnZCzyN5wL5v0o9zEduLnk0yOm
mKRw3oirpmztVOGWH2lmRT0xbd0xoD+TL5laHyuoTB2xRxT6GDYIqVM8HvYo4LjwdwO+tuiROIyv
wk/bKSpkcWyZLqZ+JWPyMC9oxb/kwIgmQBDL8EjN10lkacS5SHEwWLPUmiV94fEUcvKiIPN5yUeA
G27F9Qd5rrGAxeddChCo+LwuWhc16hgfqGW3H9fGnvPJBNrVnUummG2GPeWlSty9aPEzujPoOl1n
V9y4HVxLsPEMcDDEiy8okDQw03+SpiUJapjl4hALjhFPLi3UVLCG8S86ZGKc858bYtX7MH6xbAWE
KCrw9hcJVQ02hT0CumhHkcwTSzYbjsGm2X4VDuvriVfzfA7n5Rftv3VahmKZvij5iSBGuRQ6F77A
WcKrg7l+FuIHzDPGpOyXmZKJgAiNEvQLcIm9bkJvQkg/VvkNCUyCXrMvoRJnlzrJrhyta6y6DHCx
WelNgaJ8yb9va7pUz50SIB2rP6oW4GtpvIyQjD8k+xpjNdjiAx4BBqGEMwswHTRtPfIt9ekd8jF6
2Z7VdpXtnBh5Q42sSrd8kUpl+gD3gytiHGdbW1ZWp14Ui/HKLoXyIl3aK4/g/10WCM6vtnRfyAbK
QwACGSEE5wDv6Z8gkKR6FXgnd0t0+OqNluQQB+PEVPjcX1OV5v+O+iEdQpttuf8BAHIX1TxXJCjG
4pAy/3T6gRNCe8lnHpB2atnthEQXQGSd5iOk2mnvjKwR2xUEu3nD5genVukQbcKTqs3RTkNax0qC
gbJi1mIf8qKvdm203gcM25xf+9h/uJ1ELHZEdO8V4WrYp9rZE2gm/fEh3cUC0bduOnAAUFIZFgS4
aOgMlu/o7+7I5gjtlUldRg6jh4/2kTjbHq2DZlzxok2Hcu9Fko6xJEvwH88HazqHyzaZbMWFiduJ
/8QUpqaaTBl6tShVyotfEEDMrLMVK3Vcw+VL7t14Jo6XmoSOP/jhGznlVICD6P296Y3kQVWfvqcH
9fTVgoXzyKTn1+POL9Bm9V41E3WIhQIjJxZ7WJ+TEs8IhmAIbLXXa0bivwOVaWaUb/TRWeY+fghd
qWWUnEfBeQKljy1dmgf4F0Uylu9sXBBCnRSVDgjggVVKtoFt1nV69KNEr+u1KGZ88vIJ77CJrmwl
qpFXeL4iZNEpFPeyWuRMOeAYh6165WA6JnzO4lp+AzSwX5Iq2/UFiufLXzs8m+QUils8MKoDuTys
/hg//36rouPVLSgbTkS/5R/RE6N7GcXnBiEo6li4XEH/oGyOfkdNC6EJFVJOv0jjeWFUteQR7BCJ
i/XIKAVq7YEV+T2LR2ZjTBpIzGUzZjrx4+mblvrcjbrEZevb2WUc0V8rz8/BqerA2XaTrNnf2j0D
Xr0cLecis0J81hSVTV3EA9ocgoe7EDD0YLhRXHuPbo6NKnKnpEtV0qJOWW2e2u3OaqCe9kbeMPSV
atZNFRxwltABub1Do7YxCxsqeynd1ZknwfZS/Kes+2ZqQMU2+fGcmrpQOmm9uxZOEVAnshscfOBm
K6P63J6WhUq/ol0UeaHJnjslRvd3O7KDF9lgHsSd6mFOI53hTKZKo5voyxUbaqZt/knfSreljkZJ
HN10/bQLTixbrEqcrl49O5TR8Ky9BhrYD3+0dNZ5+r8+RqB31fhrUOhu/3mfTV0VAHQufsEUjFbu
3zZqXBs9knmxpLOyXS42RWmN2laDtLkaWNOMEwl2eyLHwXQm/DR6ZoXPKSx9wrld3Etrm3qpROZR
4VBnmbtVPvM6vLv7hSR5ZspGhu9ymtnyFWEDs7it2Nl7Nz7vNfHKPEsqpncOAnE74rY0hFjUZyyl
aC9XM6PFP3s8OsZ0Jvtfph5TNZ95sIHwM4lO2pXp7GvpFQ4AUojAD3Pxob2ELz/IYXGJxcdIE//6
lwz/h1pOnZxKGHOEYYKw9bDc3Gvig86ZgHOldMqpR3iQ3lm7AekvwFpkSQcL58CH6OvzEQm6tqGP
ytPiDG0M0LCyhKnuK3/N9jCxH+mz0DlOfQUg+X8MFmj+pzgsk5erOfqMupQ/u7GVMU4ZxeSH6aHr
4pSqPQqrIFnQbr6LR2/YwykzEPn8EioBgWJlR7dCS7V422YKcKmwrF0CbNZPtL/69IFbJNFls8gE
E1KpYaJ/N9Cc83DZoXxMgtUeevu7ySAZbZC3ixPVouXWvVc3Niv8xuvGV3MqDDbcD+HvEMEwt5BN
qM7Okb76nqKT8nmeEwvcobq4lNfmVzgr0qtOr4wNG6jDw12c8bewREz1ZB30njQYHdasb0rqqhgB
zzI3obeRLuQ+irQ5fj40ZBfpEMMvTOoK2NE4M4x0RqwfcYZMI30id74H6aR4KkhfZN55Avwn37km
qnNle3oUmCW/PhPxdP9FQ18MSF+wnjroTfu7Z0C4Bv6PO8XFTqmkwW7Y2uc6WNR9XDOF6oropj9a
p3m2h0bWR0Q1ZTqMd0tCJQiqS+b31ZNgE1fRLSq4Pm35uszJBpqZZHt/7BSSuoDUJieElJDNd8i/
VS5UbMBTPCfYS0ROiZjpU1ijlrUGvjvD4KsGV3ycLdclVFCP7SOx4hW2J9dZxsN4zgoo/iXvxLKh
OvCgrLZU2Dof3XOzGB9/X3F0b7le4l/r6w4ysu5uyumalsL5gat7dV3w9BnDecjGSq6yUGPEHjFw
Dt+L3zFFV7JAkM8AS/KYUWNcXwqtjrFqc72jt+zJTcgC+ugi3MipYRD2gE3fxCvIRvd/qrswBHwr
sCJvM1xDiF5ajepzLpaftE0hMOG3zLHDa4NQn+wfk1t9upD7IN+//U1P1yxe+QJSuuJsqOPGrPyc
Q5TkmRrz1KD+ujyNkxRajKAOhjyYml9Jl7a8nmv9ILHU8lSxxF7zZRDMNnnss5Jn7KGNogpybNwj
974XcHajBVcOYgOOkYz+DaveD7qzUQHuVdkKlBJL+1vddtcxw40kymrrpdyMupZk/vfStSn0zjCs
1PrVzwm2B1dbGv9qydBrL0+eIFT2tDigbwGY4UTdi9hnWVOM+tggs3s62MCrXpk4JHVN/QQuaZWd
f9dmUp2DfMtTHcDtPzFNnGMJ1y8d8gd73972Y3mXTirwuwamNLssGwx15a3X00yoVYIUK+0eGeX5
6PXFy8br6sqyUeHVHXupL93KWnI54fBqJjFioKl+z2VWby53inuyyCLs6k/1q2Wnf1RwIV/WWwAb
HWlX/1XxaTa9fPrSpNcUS9LoJsEkfYZinZ6eVzwqSSxGzp/GX4XelT7qFVankLOYNVZHVqg/+tfO
O7+yERzazHZFNPgdm3K8wQ/7rWjgBLBrv7bzTbtiADACnyI41mp98TqaADq2XBDi2B4DE0QrTupx
nvNnqc5EE8Tug7lJoyv6pa5nUc90Q1MQZD2n9ItWFQ/8nxwA/R+idQxfSd+fyiCXgDBuSn8CHXIp
P+BJgo7+CwKPmzMF3D6j72DMkFJisyQ1RlUtVciN/yvUSAL95ZBr/94TzYC5hwakhRJZCZutBC2S
csOLMKfAUyAmd0ndgSgGPYNIJv2yptp4cngzuFh0olbxZyGguPGJY8Yhgkbj6hRFjOXSLcXhq+yZ
jArwQGZULiplWEYVFyHi1nuNI5UFdyPhS0O/U3ZeT63CN0HXDPG64R4UkaqJ8vRDjRhBJW+13XaK
v4Jn9Zi0uBR+SwkxV5QjIEwHF16T/xnh/CONqRxD4e2gRnL4U/56OE3u69u6HaukbuUZbEwcc8j+
GbPD+ZtwV85tPdGTheFjPRx1XYP1DTgP23JNqDYHn33bfh/3oAh/J5BjhiIOXeHboV/Y+N/oLsIo
441TkZ/MRJIz/deZmaMCBex+laloJQuffWv8e6xb9sO8DoTTVKMbHL0NsNG9814tUo+QuRBMENLX
QkcGexfLWAgtnjH6bxWXadGdktauT40/5KoMkuf+6Rw8/yeQo/tQ7iKUCGzLZ17WqGh/pCSwNt65
TMJ2EpcwKpJBaCj5sLUFBNVq+9uGEOj8mw8fK13GSbkJrecrOVKQWePdc2XfiVTObFzIwXbMGU5Z
hpMnsnju/VEEWHLvfPwD24iJQrK51VguMjItLbmq3hRVDgcQx3JT7rgkhMFVoOdq0KPZNGHwMCtZ
CraRGL4U6XyCqU8cXAKDqDZmRZQkZAfcrsy5y+qzvxbmTdEKIAHpetIiQMOrT+6AhnZ9n7Bhybax
Rw5cR08UGqJAEZ8RgZ9eGdBqgl2kZmEO08+wlbvLHzLSBhtfYwWtCfdv81KxY6mcAQc60OFBpk8q
6ez3J/9Q2LUMCC0WPikskbT7XqEQlP2ABrjkwRBSFfSlToQg1tfqn1EGCjb70AtZ0rFJNhpcaLSm
kmlOb13CItTe4UbGhwqLB5bXk80oKpKS28YQRbrjz2kMcHRDuiyvn0LYgw9xAkZWA1mmUnJqqsWq
0zYhdxZN3tG+mvnr0F8wygUybnJTb9s0R2fwxEEWbIAv0fMlWOmQW5g+wGmFXLw3XEDtdXAEghCt
ThbUKDovZOBrty3pWhIVs6LNjwIusBMAPXX6VtVGzTKLpk/vdxMTpBQp3ZoUxM5gygCC43rAZCtT
A8u2dBleHoqA+YLDV6iUCdEuVk0TRHDONHmMg+FzYitto4QtYOU0Iwiwae/9FT9Lv6qcxgfrmrGI
UkPSwmsQ1+/Mo0bw/yjSmyVM7qw14AliDX2Gnoy+KDvh3iRJZKEcmz407OLfrdKWczoYw4/Nr3eK
7vphdj+A+1UVF2vnyXTZcaPsBaMSz6r1GDCgKijX8z/GuyHgTflv58NkYtGhTq6AY3P2FuJsFNmZ
oZ4WZM4kp6+UVf4iM2bez9IvdGtcv8l7vC19Ry+8/CnoF8r4QdZBLVLhs79WlJ8JAbIs1xZD8efw
413L1+6RaJ5cD67It7J4Zj6uYU9fe/0QIUG69BELcHw62vF0XUmE4ROzwzmNqnfpWzuDE8OhCR5p
w27QRxuGNT6cWgnsRpQK8IfiersKwODnPuDDklEuddmDrmoojEPfhtR0xJfCRHH2+45No9sE4UVt
XDU29M5YZeitwqBs5BVEfhNnZIYkMYiYEA9dnIZWet0joV45aUKS22FgHjlYoXe2i7P56PhdDInT
F5jV2AL1cHiYbSLCPgLOpCWmS0QOxh1Dm5KLD73yQnzXpImPXCGJ9WrLUT0i87rX3RYHBf7qkFzG
AvKICC5nPDlwKQJiwIHxnADcT0kuQzq0lVE6UK9MBBpzWGJ5da76LdkKI9KqDnYeNMz+k5XuUvDo
9ZXFWwDZ+3kxa70jocTm1qSSJ04aNJdaZ3hd0oCZHnw4DCagBgFxJ+Y5M/ulTf1NJKTOTSHXH7/I
EjeYkP3IN1R3xfYfoDBw87dLlvMtBrM2tgxow5cWRpW/J12p/22I0Nb2eENUNBOlDWNLAL/NJ9nw
uaqkK1LVI71xXDJB8sthxvXETu5TkeLA9yyq99fNWwHHKKo1CGKgN3Yxrv7Ksxag6lLcJJG1/ac9
hKAh7SL7gw5jqX9UXxC9jseWSSWIywq5iuNuNzcdPrkKAm41TECW0hptXBl9pDEyOYCNCrLq1UJ4
gagpLdjCsNeC8m8A6HvVxsK1t046F0ecp1lMb0m4ztwWR4bwA47eBGjkxGrAwLjdfbxUap/I5RR+
/2cTp4fQaU92OszmqEfU/O7yL9OCBDSWYDGSSPmMmLabH9NOOrXfo47RHOcnFLPxQDAJ9yPT4EpG
srmyxFeGlbj92p9jcXC05O4rkCqeUgVnHhNOo3A13HCEbEAn8+MhNrC0KfHngA6SZI9XveYg8XE9
7K2+wQvJn4U0d3peFtGnHv9dAYv8XkAUeCJHo/dgXxd82prpbdJm4QIbPnYr7hOrRKuzig8TqoJm
tU1r5XLxqeYKBWEa4U6F84H39ldOVgMpP5AJVzGYX8ykRa1cS8FPpuedervUzk4HJIffhwOpybIV
6gTZIZTkb96B97PqZIDgTD9vxrwc50YWTyvBmhnnQWejSGILmQzfqInBQ7OjGgQ7LJ+DBPbjAfmk
MmIqebSSfKluKRdGpoF1KPHHrX2cwMtpjNJP5oEbzjEW9bxHOqvJT6SCSVJZILLDPPgYnqEtb9id
IHpU2lgar9xY1EJeIa9B9BVAIMKKHLgDihv9QbCzmXuCg/MSWhtrGKydrjVtPaZHqx2+owS3MpWY
Rclv/w7CTvgyWBbFu+VSqt07i3C+B38Vq3c+THQWM8mX6hOU87oNMBUNwRg6L8+uOgSuTpGGyyyW
pTv05wDW9IJP9DHpWIG1LrBNu1hcYqAuaz0AgpFPgJTfaZv6hjVLcZJnJGuMQ1qDNveyT9442enM
zJauqXzrJfnKd9l1ry7T24CGH2rh01J3RF9X/ws5760T+SH1F/tbdWr5HEfhD4q/2WAVR3Sx+1Nd
fsnKeEBKgGcGY4ctHspEiluy4Lh03/ef3vuv/D7do7CA7HW6Gln+MkX6hi5OGAztk8aEhIwFe8Sv
fZTI3UhpZOJxsSQdnjQmEpg0YKFqyYnkicdY7dl7ITymh5BP0jezwyeigH6FNQQsJtwOeRNZsKLy
fLv9It6QfifVEVgokoMmtQbQNqyBThpTEmp9FFe+BZuV2vKsENNRjptWLRUboUWbHZ3uUqlSuSrO
94Gtr1y8Usvf3g5O1NZa+IhOY1yWWFE37DJoodR4/ufiUzJG0jc6q6sjb0k4FmH+wNqL7hv4pt4P
o/0rKCWteDuxT1DvYBS3etaNZD6ECN1OBUnrBdN68VOoWBq5GbE6Scfm2jbjhJStgpaEhxbjA3VN
NpFKoQto/C3dpqlGzp7GLkzsv6JwggOyBMVJjI36UO+4Cn8eXrIeDcV5NHVX1JpTkkzUGRXFivmU
6aCagOV4TnugGNgVkBsVJihFvYUl0L0GuhfUiD3gAVM/nLBkwMwENrkmk5Ng/dHYP8htLrMJn/mq
aiG4ESaGzbZ3KsjylcKnVyKkQpO3zjLoto6iJUAUMTdmlRUlFQyP0+WFdOwAggum5VR5d9ID2CI/
dqvTs0ASaIlhEIfv+NjAwUiDLpzryWoIkAZtfAyqfcNf2IENyg3gQ/x0f3s8agqTfsBzzEDqA57Q
AfmHOrqA1E6wx72M8mgF4DB84smKBkYGEHTvUOi7X/eBTJaeA4WEdRCSu2WeUo6SZmZSIYhj4diq
43Jtpw9FnFdX5TNp66Fh/3ryvOiquPYirQgn7pcQ5/cO67F4BHeg4RUiN7A/CVXB8Ko35uGPl0mP
Eun0zOK+SbyLIrVq5VQSzp5BT0PUmmZ0N3kYv35Bj8X+DJIwNiC3xNsVC1nVXBBSFiZvLyqarCmh
tXh44vTil8R8OyLzzu+sYP8uuFo1O9oI8461TfF9m1ZJTCpjxDSyPo9b7C8Z/rUcHdiQ1XFrKsMX
sb1r0iRNgcbYgYU7JcU6Xiuke5KL2HIkLYie33PWyLzvyN20WJzE2sZQyu9J0NchvrC4oZy4vRHt
HWUE8gLzDmJTXybVB35aSIUz7FnM2cv4GwJ+J8NxgmPlBhifmteyv4+iwf7ERHpV0lIgOga4DoiY
TmthbP/Hz3/QBqZGRy5x8n93s1zFNaOLqbkyu8nohtSQYYz7yqX6bZ2mjHh31jgyNQGaoFtHKTB9
UOCIXOLCxYR66BYgayE+1EcgTigcYENakxnvdo258Vs3TzwHmsvMZItY8r38zi4tYmGFhjqOSnlt
w1ftXR4yS7v1WgWWcQkBjnKJWKQZXbt2A5BObAiaVdYAWpSJ6979YqkkzMyIMECBy66klei1fINe
V2+dCej28yfI/CkDjgab1ygLqM4EUczkzx/71kZpe/H8w0VyXRAxa3qyjR63I0VvbPdpNqLpSB1X
qypptkiDXvQdX4gcUVe5nDv6Cd6uIVJRGpAdD0CGNMP2h2BeQFYqJcs7SwCwgFdszKkkWdE6eelT
qRJA8VmTaSEo5cN/jb/+Q+k9RqL/6E9D6R9cpGn/2Max5UpUsSZsndZ0lMLRTJ8B48llwOwsHw4j
T+aOYg0EpGz+v8CdJcgMtug5UyzJ7BOadCLb6Zk6jaqyytHVWhEEwzaHgohcxHpxy1fE9ExD+Ipi
8Pdoz4X5JnMh/t7GXeU+ajgNT0XodxpEkhsHJVer/aHJQMJi9sHPVgrySMWFvu1YC6ljyCNkprW/
UTp0aHxpDGh4ZHmkzilaokl3BfAzTw762PPA+d1DV2Go7/uxVSk7JYcM8BnuuKiWnAqyhkdV+TMq
Hax/5WZdFd3u/yFAq1txz9OYwEwxsaP+cogjpkboE5rZ1zKrgaBNvNqVjry3SUDgAjbXi3PL8skr
KXqdJSboRFa2024vTPGMBMob/3F1QIs8ORV8VJhJN1481lZHKDXDAFcT2iNMJkC2Ds37DUb/xray
/zFmkzCp8zjnAVc7hGot3c72knnCZVcYyJNwUG1apsko+lypZkqUhdzyzKimrN1Z/mH4LzldZVH+
UgxwTgxNBlBmW/M57EyBKH7kbKQqN9NO+tQk5Xi8J1LpAUjg6dk+ezxl44/et7ttL7fbyvWf/2tQ
E7Eb1UKJys4TVClXNSRXetSNZ1beuKLWq4q46fAAppAdyGcl5ONm4z/mBx8qyWpWPWMXg18PAaBX
tuh4MvoOaKE4yV5o0RHRaSm4Lgc4JfRsh/Hjpwbh+tXS52yTbw+/iQhiYFJ4UHb56poH+4+lTl8q
mYEtlm8/UZnwkFnRwWjGS9VkfktyWo7S8TOqCg5tJano5D+j9vDzffP+u1ZS+TX9wRKFyNPzpVrV
foXpceC1d5waE0RvtOokP2DKOb6OpJgPu/kL/FlaIzq0zBBbGpA5Y4QDxgJf14ZVyNdg6FDx13Fl
S+38SfUDll9vRplqO6iUH4oU6gqg//XVBtE4khrnV74D4JKb2grl5+RRb0i5k2Z37VHkYG8WSyp2
0Zj7DOg7NSKuZrx6Sft9eEi1rV08TTNKIr1a89Ff+UZmXExMdcil9NaArDtdHapFty/SfUTSNpgJ
HUe5GN5DMPGudlTM/TWRaU5Km3JJgTby0d2h355MOGU13jyXJldFIWmYlLKdBWJ7q5enk9j6Y6er
qdZ04u+Gln0IFsChqimlsFRBqfuQEYpn/sLAEVp1sOVvARWP9J8LkWs5zLs7LvaXe+G4Pe6bysZJ
UDIn5+MTtSqslFUgDcFdH+BwJRaU1ebndhZzTyDfSzkdxf3m+I2WG+imWIkHk/y2vfJRiyIfMp4n
ZWDqyj4hiAbGzkhr9HWH+Ff47zR1b1KrK7e+gp2ExkOOBazzwB6z+mOF3d+6crDAWUpg7HABTyHQ
ISRzfAsB/I0D8QKoaVb+7VfiTu+evMMnfJHesWmCeeeiY3530jBcqcYUYN2+lUMdUbm+IS5mHNUw
6iZR3VN4PJCc05MFgqOJIdDQw5JMKXiB8Z1oZTXjQnF70jg9JeQodU2bKFJujQoGtaZUDSAyZJIh
x2XMKOcjdpMy0X9ADtHkEkKT+JoDjf2pcfBTgSZEZMci7TR24n+ZW6DerTQzNgxfMvDWNr8BxCYc
dH65YVOgeH6wAjJIu7x4HiF77tvzE29hj8hQopL2n88QorCYyGbSAULu/aXe9Sji+VcfBS9N69E3
FheXforNIv0seaW6ueTHmiXs+LSBM1iUVpdVOfYNE708pmGD9s0ZF4Bqj9BnimHRopuQqhGaCEZB
TCloNec06SBZj8KiyRWD9SvN4deh5eTqT6ls9gj71PbMSvyOtqvdqXdJ3QzsRPOV/KUR44ORQHM3
CbrNKP1VdbSEs7V9Xn+a8SUky8H9bTwBZcGvWl1P570kr7D9c+O7sZdzkug0Bw3sCdFVNEEi8Y2M
tPbtTEwN/mILq0bwbAVVVDFwUhJX6dLcJ7Mjg7x6gkDQmIrlwhQUtdtvilpzCB7/JizygjU5Xyzx
A4vCWcTyiMOiA8RQHYkPp1ValDmVRaHyxy8BDN9Whcpv0V/1WTdVrU6dc4BWQXDEv2ClH9wiJtgS
xhHjUqniNxAuGqJzm8CR76L8YDi/tNubWrXZJgkSNtSGoVTVM1MPdUk/Ks8KSa3EYRQUQO3Yfwj4
T+OlmN7EkWGasFvv4+Cz6gR10O+J+u5kQ0q8g+yRZVibEpf8PTcThW2STVq8ByiXpK7mujq0AS3+
gKlAvGUJUmukktTx44uykhVd+f4HV2vxd62qiLvp6P7bWi7hUmg8G8Qp8lL+D/GsadZI/gm1260d
3x+v2ouq+4O6X/TwUJhRQt0LZDsbORXxtC2HbKx+QKDmu6Xua5I8Awvw+wKtlsgZmYN9JY5UjEan
LILb3RHmqfUB0mIHegN6Oi3QlBOTYCXk+dDwwDNvBhykTd4LL/ejlOCirRPzoWjaRfZX7WRevHjw
dqOXX5A6XMOt/xtz/bzMRAxwLcuUlnjb8d37Ix3TMDGBfjOkhRDXjtck5HUuoHGtlLp4Mrw4P3/Q
ZQXdz+u4A4BsEixt2NmnsBsVVYnpKrm3NisFe6/4YsasgGQP9cBqfdSGMhoIFfXPs0j3XuevQOxW
m8Lex6dHMBCtW3FDzuQWD32NGW63Ju5+Owag3yyA2AssfRKRPRiWyykTk8f+dB77es4EVNlJq1/I
2UIb6TELlh2XkpxgdDAv7oYluEBIO1+iebl0Twb+YpUT/VUcKL6XJiLiNo146DZ5Siyh1BXjyp2T
/EpsmwppbPqsCnAOJPyWWa8MqR9qKAlqz+VNQBN+g+fdB3Tg/AD0GyhGA5ll04ZmGvNr7Cr+XWoi
4L3fV72Urnxr2XAvbpYYZhbgrQPqATqmk5qxj45TX3+obNa+PDGPWwAeOJW7DvPQL8/wrwGpOntl
kTAgVFo2mtSwJ8NX1sX/IVMk4n5F408qB4eA+IxgJuCivPn9S73vG3lo3iXEbubjkJKes7eCVYEN
T8jS8l00swiGC6ULVJdgaiEJ9AQO5DilpNpkEq/rp9FODjRI+AzeQRNHi4+XkM7OMbPO6sBsCdD0
mQ11vvSJuyHLNgWxyw/ZheZzzya3DpgByQ61UP4SETa1goz5N73WWUjsTk+4a04xlA9iecV1nQ5w
co8Or2hZ5Q6Xov4yqFNkyOonG4TF/V9Lc3T9+CNoUnxQGTTQF++Ybto2h4RAEuJF3GHjYoxu3sza
PCn51fjzIWL9NuMUgy9Ei8H0HNGgBpi9/qP0PLW3EA9lpdN7H/RYDTb0sI1y7iKwUBFXXVLtr2GU
t+zUQbcDdmbZxd5/q0HF9bF8KPpuvIm3D4rq8FWCbkCg1gq9D2SRkH6rFgjQm6RmaJVeWFx5AZTa
44nHe5au47/Gld82RrLj0ssE3fHERYoFhm3M1iK+LbvC2d7Qozy0MnbrmIkrBW7PwUeVKWUzYkFO
nkUlzGD1nmvhoTtvSE0a063P7Fz8zMDRSzuiRJxFd2GLO+ikQDuyNmgKAjEanN+5qM3ySWv3oRMQ
keGoFDCcQ+NznCD+EGaggctGHse12gFJc7l6BH8KuVj4uQaKcgj3gWfzIbPZY1+iq8R01blxwyRY
VgGbNuhixCgTC8uYdpQ+jcPvGEFOr0jhH2ZXtP3bPk7I4eO0OrKbAqnc5pdScJDHWX0TQ6hRiV7u
OKFfE6DzXdRqaHGwxFaJV7mA9nmyNyhu0hXskEHP4tJPDD2KocjVr3Q21OxZZMV9s6fYarP6kDWN
+JtLoLpy07XovSUmgpcP3y/qpz5cQ4ocBQ+Kk9GSoSvwK6G6A/GSPOiimqpoAAqKDChJAdXfE1DN
7OaEvD5dTFkJCGHhuysMGVG//5btQ/u8+WEskrrN1XyMDH+GxIidQP/ZizkW8XZp6lRs+QzK1xds
99PC4ao8Bu8IUje9m0mA3S3DRzrSczDTX6SUB3WjjdL8C2fK474QKEtNDZsUpcrCHnlquF9igCmv
Q88TU/1gZmWk0AIDM5qjpkAr+czQj5hUV2u57epKCVPXdrKMsVaJeDuvQZxmDA+mZ1XWBQ59q4a9
ALmCqPKsOHAyO+trdHEt0EEE7rLQVzNBu1XtyGjZRKHPKR9/Zy7Vphk7sh7W16cycxjh3AEKhLq+
WMbIwZfME2hgcz+aH+8hgvgN258eItKvqOC29uavOVy9tbDq+N0oXWxBRCrVPCxUsU1qbsX8lSqe
mcH3+GY+OvO06zJ0h1p3wujgDa4w9kxCvRu/iBAqyfq0gz5OjCuPnv8T/ftkQO0T6Vuyv+0DI0zq
NjAw0ze2Ot9jyZ1PHkoSGdWdEuBqHUQs8lI9dlbEsyJ+uK+6f524eZMlhaFiKYBN/BH1aBuVfYov
oIWcgk0WCqPgMGc1105l3Fpu6z5401A9HKV1691ongnlAr8RrX5Udr5kiyDXwn0bzdsTMepcEefm
orMA3Vk+PRnMiwX9vTrKEld3a0gX5ev0TI+BBDsdHFTt5+U+YUGFnDnIjmkj9vLbvIhWg8QhGd0c
mG0AYtf7ctrSyaQ2c9FnTO5ZAQKjEHQi3wdfIaCO11dxWmCYMMqqVa4EwlUZiLEHCzWaiIpDikus
yeGDGbM8ovp3qX50/ebKr+IoOrM8v2TXSIAd5jfwhcf0Uq5MOR/ib3ikssPN5WEfwUoyVCsXTTKE
lNhNccWkVigD/i6UWRs6JZccxQLM8mRmObGz+znNM5jUK9zxac82DGkru4t3mUFDzBD0jfRBJpVv
JhMGjHksXmpDbcyKPXY00DLpPvcVEhIQm+KYG1oqs7UDanp1KMP8k6x8tZ1mCfpryp6bvk60n1XL
uNT1N8etDmwA45mrD/Wk6dWHpLiFgLxrxBsZQwRjm5b7fGmp1z7p3HsmtkqNMIj9SGfSfFKL1ofj
dnw7rkkv5dHiVj+4wkkkw+a/hOdtnkkUMwc9GwgYqCD+VUTrr9F/sP+WXwcQoLoD1vu/tSBT9FCh
mhoXVwfZM8svb2IhVh9KUwRxIvRUcyV5PS1MBVxydJjGq/yw5l/jIAZsIi1+8zQmbXGiK8EjafmQ
gTCTbf+4PQqrN2gf4epH5o2ermkBBY+NPhwrAvt74B9EnsVyNT7jCNHCQNHx+OdKsyM/1Byw258o
119dsEDX/jAkvJqcvvEtVvCdsMhqslcRyy7jZDe7XA1iNY+Q17OIhTPCqgqqhzX3bKmej5F95v3w
ASQubfImg4GmgFnMODdTPUItpYrUfTL5esGVZxxG6VEhdp5jH6bQSsQjqZU51+MbZ9ekSjamJnK+
74AsF+7SKFl1gcZgLV6s+1SFQ5x/HeOo4AgcuexJimX0yZZ4F7K19vB/a7dVTZJbwkoZTvw6VVNu
Wm3R9spZJN/DY7ycISh4rZWs5YrnZxT6tAiGLkkc7fqXSpcnYD0ImFr5i4pYOex4HlszLWiQcQP3
dbdxOnITcOZW6mUe2/onCCEwnHxHTqMoMKWelx9lu1JQWAartXkG0IuvAmzgZ9/XvAj2lhdg5bYD
MdpJvUO4olDRxoMFyVDR5BrvkyUMG60rD1itF49FkDNzdct1FT8CD2H1qapyMsLfytVZ5G34vEsg
xXQmS346uTRg34C0Ma1cJ/D4FDZoNw/pp897ygzfa/15mmnB661ynlxQxpsqSX7AcmcLqqZjZ7Mm
M4Z5gP5KU7QgSCIU5BNxhBcEyRZEhszobzhTeLhXqjgzHxAIl2DrkWTJ4lDSvvqqxX/w/YrDtBy/
BNcd5DrretuD4PsPzxTG5hIvrTSpCaxuG4ROTAxUYA9uC0GKm0IXVNE2I2KgiOKXgi097chZLbOs
XDDJvCeN6/SxrCdkU+3PeZTb/XdCA0BpjVAUFCoRZRxO3aTF7Y9ZwG2YXDcZ1LpINUYhQyJbM5Ua
LyHs0IZsEi7B+PzIJbFVENoaufFbVUYhG499gDmF5nMRFE5wk86OHU7nT2A2Lf2vhndZBr+aUqhY
zv5Gi03BiF71zZZvse98Uwh+qKgSANDXqiFDV0W6rZQrhTLB7sDn6wZxlbiuY+ReXSLz9TuFZTDD
3zfA5CXstFeYzEEjsyj2s/s1PehFtc0z7532WlLig/FkJs63MiRbN6+wBe/58Hhd588nxrVyZ2bh
oDsYCw+VS5czfqCW5EhAJxUbuiqgfLeEyS1e3Xj0G1LG6cK6AdxgQLIQ1zKytf3wG36yOSoyCvuW
hP+nXX0e3zaLOCp4qC9UELn9gRYTMuO/tCuGYOsGCGlDd/ADIzt/3wnS4avOePUzAzTvW6wwcNIB
7nXHijx3LVQvx98AEVLXF5T4v4dBpU2X529FyngY22/B+2u9uPY6eKjN0z+REO1m3BApqY6/83KN
qfEOMjx5MgD8w/yPHFkGhaDaAE+aOnXBU6zJwrDDANEYJkevXPLzlGYRCA1rP9jx/GmvFuQQcOm9
3bvz47yg0YOm+yYLCvL0xpCV8paiWvCXG4lc2wv9bBe9V10vAd34sU4aP/9/xudw47HtXJehiqX3
NnQr8BoQf+G16lEgwaEc2soCihtZSATMkf2XMGimIxe+OvkQGzT+9lk3tZAVwCbsQAVZjM1aBulz
YDD9FhzZcaRQ6+uyH0HHtbAtRETj34+kfk5b2mMClHKoEHAcV3Pvy/3XNdeFz6Fxarj12stswOIX
OvjJiRBeN6QqhaKe2trM/lng3PFm72NENs1DF+V/N632+gY/sQPCRuO017U40zUQ3bfCOTuYeK/s
w0abtE66gg6ao5tAq0DYvy9bt7d1CRm0eJaqYCdgdN520eQE0EwuxPiiLZOl/eSg18dwxpJRul6s
gndXofOF+FiJZrHHeG9two6lVlFiPaMnmk0vA6xglyVQmzBIAIcP+JHjPGNzAy/gHurZX4CYfktB
ChSr/sJ16cpr8ayyVBf0mVYzTnhLqsyazlnrp8OZCNG+69yUktQoZOTFoa3rSq1nA3RKAMQpA911
YS9EDpp/eeq/bqN18OUWswOgnJnUNIHy0papP3NVeEgj7/qZDJ7NGXv88Rmcsh7ud3LE/hzgUzLY
LIEh6Ml9F5/tWqSnXXr9F30BXvQpxlHfwZ+XUxtU4eQSammWxSrzsf1q8UgwlOdF4AMC2FXSudwH
cZ5JZNYgKuGtjcdO4N91ssDU1fX7+TOQzkwT97w72yJBLCUoiRzvHL4mfCuUwhbrcYcpcwVNw+YL
LtF37hC8/gHhKGEuPvfQVzya6WB24GVEywubpiveN8t6ydypHpEn/EHfriAwf8EcS1dv26xXTzSh
Qgr7a+dW93Clwq1ETkV7h8kjVhUCkb3EPdAQssvL7PERJxH48iJFxhL4JO7/zn7E+e+HlUbWzbmR
5S/zRubDcUVKN/nQVkQNJWqhDVlll9Vus64v14N8Cil2ha5qRXe/Z85faGJu7ZzqTI1w0JypnNpu
mwS2uZPBqLo3fSDy3Bt3Fo1Ij+qnIlwSDqN0DPfRRrRZ4rHcJIEcJjlcw0WdxrQsikSBj9wkXf1K
6cprH55KTelojhxhFtQp0hyyAfu3mvml1iD6JpC8naEf5i/oU4U7fAlIgRWAuD134i2iWhLYTkUl
fEJc2lEpCVGi8jnP/2vTgYVG0xHyo8h0zcQZPJMOJvriLQrx5mTi1mXYK6vjTohn3Isyh6Z83/s0
j84hhfKvMshtWMXMQ+ApUhDh0+VdErXbEWs8xorZYM24H3wclH8MaZNR93s5+1QfNITWoh5a/8Qi
gs4vN75IXeZnctMa8q07aN6wh5NMsoctxBkQ6PPrPATPaortMumb/Z9NPwbmUanrAkjV9GGmjKOs
QHYshUNhsALt7u9vw01tpCNLBcYHdhR6tkdSej1biE/3ffB0NOHH/6VmZOjHvmo3L8JgXlTDG6PE
Ikr2koB0aWcPEx8tSRIzWmJmK+kro580I7eoKXrH9PfsEcDd/9ZARr2soFBGcokNukvv/9Dr8CBH
rzZvvQTwIQnqtCWEYv3/BLuVWMfzwqDDm45pndfJhUJ9MEmuz4ftXW4bpRbNGfB+dUY2MZ2Ib+7W
qdWqKXD8j0bbt22V/4gYV/PFIV2KDjED36nj0RuGmsz4xRSGDoLyqSP5eCJCJE8AFC/EpnP/+RRj
G1idIpm2FXML9kBBjlGnwvepxP0YDjhZ2Xu7k5g02rfM22t6wxParyZsEMjZC+cd5srwzTUyhaT/
X/X/Emxry8vwaLvZ5dWVQMxJznFfKwm7F192bu9aqOIEHRWzbTKDR2iBcVT7145Vn1mLcUcimugN
2MszUqtT9zbDGlHu1q9t8R4RlZ1m/YGJBHLY8YmtEgs68M3zlgGDr4/XgtBlIHzQewMUrHFhNhAH
0cjtgKeelnZ+JqUBVwlwpsFyKpLOqGey11xpbilo8ilFOskJXRUdd7kx1hiaMh3ePBV4gcZmzMR1
eYieSfwc0TdHaHxQe1Tit9VAxydMshhnhMJ0ACXwFKcO7Ulr8BPZ9eNAhFreyRHWEOALeehW1Mi/
iB8wN6po2gxXJtobVPeCCqD0okhzu7yMiljOZPJy/eiuLCGixdJfSYo2ZNMq7mlUBMmXTiFFOiG4
jtptISHLjRZhB53YdrUHp3jPdQ2/yrwu1AFpnFmnwcvt5mFZjZdI3N5y+dtvUE5eDe52c8GSkZAn
JRVma3JmRW3cHozrKNXDyNO3Wzmc+gFRhxxFhWlE4Gi2n9ZG9v2/X0AUq4VzoOeXjrLZNbewvIPa
AT3TOcSm2ypg3ClHSwnxhj1LWSDUeeN9xjcLmRtSER5xBBMEoUk2c0m8Fby2VutNVaQ1ZTPP8ivS
JakLfxP6IzzOdiaQ3X3XJvO+LRfgfJ373Uj058hChTIR/ht5C/cubMsgFxQhD1u9hye88/X3aj4j
yB7UwlMFf8kGYjFbvQUbLFyZlPH0pXHOwr20I8WGriqUkkzVyC14AcmDl8GaQslVvJyQgaHBqt9K
ELwD+SlcZ/b+jnhGTPrN5O1DXUlWT2SbQ2uijNWO48v/9j+yh7JDuJ6EsW7oeMNQluW6lL/CwS4h
9nOYUqmg+/9SSWRoVLEshkaDIW5Ko1r8fHy4Pm7QU4pNQTRa2GDFT+VffFDPqvee/ZuOpthbR8KO
SIHCL/kORETDyrcTMVCkiutUW24DaFBgcOBVMj9RkkmOxxwKbvHcpGAAK7EuLR/GpRpjalIjbbwe
IiYamny/RjIWAwcy2MfVOST7XeMPqkZVa4cSYUNxpHFQeM7gTbMstghfHocSO8m75SfW4IKKHWbX
bTmcuOKM2DVqHA/HL1K7GYwQg1PsuYzZBM61gpBJjb5AjwRtwJrms9EVh8b65yhiXPi+QxLwvFTw
cRwI0eTIhcENBsqNPOAkBwn0VRFKtHHQTMvZ7j1PtibfzM9kYx/jnKP50VXBC8DTViEq3BiigEKx
xBysZ4D97h9JrkXJ19tKlH4N+kUL69dp0bY0v/4T3ebmsrgThFvFPm8w7Y35GLHE7q46XVORzpqn
Jslu/GbHBmwsxaz2miyPgXKgDSNi3l0OWTjSacFOTucwkOI8iAfwvziZwifkcKw5pqQT/HarkVDR
E/BRv0DjXf2n5JJ+e5byGQnCnAS9Px+gKsj9t+MNm4R4dK/KYwoZQwZseWy+WBsOIghm+DrOkvy3
dvsndRh5G5nqbpNXMF7ZVpJLgsR1fA7Cjw3tlERLjeUVdZsrMX8KPDcjNEOBNYqbkZbYpRrzOTYL
NQiJEZ/Y8SbjzyEajMsXW1zKIaHavl2bDN7ZeskJUQ9jMZl+bQVGKCgB34cwXwFTzrSpruTpm+5O
xjuo4vO30e/ZKxKGibiuuRy8tETAFYlOdduLPVxfCZW7eRMZJIJNlO8Xz1Ue1CnYlDedCOKRpNTf
EALYXl5UYUEyBo2TQ6gYFcJboDxnHiiHdjeQulNqTRS8tyG4ocpwAt66W6NpyrTVK2J6JIk167Zk
1dWRlUTgdJi7EYYr9lmvgUgMTk6hFF7Aezg61M2BtnxtPGJZerrwtpoR0w2d5/y42VTJH7kXjX2n
cFX0c+iu6FdltLlJc2yh/a5MsQA5jdHPAzfroWwFMw/swUCVOgyjTXmL09c6IE2LhIFsVwDYUYar
s2tRlkf/lQ4uiDZWJo+H/LNYvsmoyKE3u0E2OddDVY15FU9K9r4lRtimRaItvBvFXOuroB7Itjc7
ifl5gbAowexX8nM8bupHyWcv6w9/2MaCAxyDemn2quTVnaB2QL32tbgWNETdPFQrN3pchd9UmD4f
o3frbeseyOexWP8omC1D/QQzAwDVqAKwoF6Wgm+WMd4ES3xHd47wiruJbLoNhf2IdaJQFgzsLPIc
w+KoZOOK1JOkyqal6t53wDMHwSDMbnO6s+lvQSlI7ipWbrS4wcnt4cxv9l5f/dbGp+M1hy8isXeY
KwCq8c1Ynn6J/2YIfIBaBx4XJO34KLVUxvOnLAZPR3aDnn8XHO4JyO2CzOXDVcvhl8cAVb8Wq5Ov
2kPgNhtPCVMO9blUTZWQVfav0T2a7rJgLx+ludn1SDwmqNhFyF1r74TFzUzscDIhGR/TxcZMrDrB
vPFurUdKSWs5KkUUDhJ1ZQ06dqJfoEJtINr4io6DI7MuLt7QEwKJH7KD7ceI0k7P85nFzW5lUheR
kyPFTZgkNG4FMK/odbtPiZo5iBTLkRFbsj6mYo5fOFpoXL8CaWgQixwwe4Sw+VRQKwtoYR5sufCs
sNkIYy7o8rS+nTDMePwFtZVTuadTy/POThGwfgCn/rdff9u/W3D77/vRmbfFvmBzIFKX11KojbVe
uD8Rfxn0l9vkAixJqOFfJICObJHtkGfpjTB45307nJq5NXt1+0G5Cu18zeqpibUXOBiOdF8F3awr
AYd9ZZGknMEuXXYSF4lDb5Um1J0t2Kcx63zK72S1I5Hi8N0RssiVA1SWU5bR9dw4y19v79Ccg3V4
oAR/EUpXLK8aD+AlBwxXx3bVhnb7j+QnmuSbOVt26oc/D9bjTcYoR1ph9mjkGc6jQgv0JTSRc+wY
1kPPh3o3U3sjnff//RxgvkDpjAFIUOH64RhVdLTbMHBi8Zw2pcGpwlcZtaorgJBRN8xP4FpjlcLF
IoE80FjTv1g5IixRuUwH/f5XxF+DwT6aOtGKK4LMIQYxEZB6FNoAQIHqDadfPh8PYs9um59PnFHN
7nBfFNKn92sK/KS5RHqTeQ404nxgM6HBJRwXYH8DPR4Rv1pF95Dv3pxdiZAneCZvav6JvrZCcPC8
SneijJEDO0IdNfs1xq4LoKlcgNqU5j461rm1QGqapTkWyQ0yActWfbQtEtBYM6brOUVrYc6TcCdK
eha3JuJhS+KXaxO6B6A5gb/Lbloyb6g3YmhWiQ13V38WwDPKS7FQtnZ8d6uRwIyLIneeT7Tjnk8S
6czRmADGCLJj8lcOUl7l/1jgZD5L1I3nnsYDM7Lu3xT8IZ/h6di9JsOcPwWk1WFueY5UJn1QWWEz
kJF8yWdaSPbZWRYuLY8aU+5RQGp6fi9G8j8zpMM8e6H+CuaRynRzxlYDVTg0SjnpFLE43ke7pYk0
D9UeNzYVqqmrQv1GVMh4ReQsH9tNj5bg+5Msvhu2jo8IiFHeA1IHJX6ocmV4iApmmBGhwiT5D+7b
8fD/ZZTk80oSJktPEKAHxSgswQ0bws3fbBCvGBM7/mMrYAY+pXAgLv1bF5yY04eWKLaXtzBUC87L
c5lfZsksC+3A8MD0htr6wgElNkEz8kPOcn21L5O8Xcz4Ih0PLmF9W24Ka8lPA1rQtN2u7V/kVIZM
M8sqepaB20OWAqqgo5kDHq1+3IC7j82odc/891RR/7SW7eFeg1k5zcr4OBbZCT3Evbc+noe6Xhzp
rW1NI/7BjJk+6YToxivXsz8Px7EshyHt/gIVzdzfK1vwsxEvmDwMHNOHCxLF2zDE3OF34gIQci05
/CzP9CyYygeT77JY19LMkbsotkXFA6j7vA1F5y/JKZSLEEnj27fWNpw7KX6dWDk98xMmT6xZ+gPe
FyIbxHfTMUWK9SCb+YlMRqLf/o25D2uw+UEqLXuOpjhMSGdgy+OUqjNNLVZPwVkLAoFLPUyUuqAG
gC671/cGQroltTHn2R2HziewF0uRbc8CHpbjUdpY2S5HeimgeXqAfqO3brHpi+2W4/DZ9Gd7ZMMz
SrykgrTtYVnV0/Wpx6TVdDJBaDr7HIiojdkSmcLhInEql7TgjY0Pj5aOsXRRDeDmDbD6BhcDxrAt
bjvnPp7sEExp3lirOEXn6Iw63tujwgCJkzdGCXMPK8bzK0JyQVafaa/wLzq7lmQLNRGR/zscyrsI
6/TWH27OUxXvzwMgLiJWjXjOSyryAHrOD7F/rGm6meBtWqF1+LIWOqtX4U49VlyLm9eMD8Hf4oP0
AruVvTLWIEAhBXu11lm1MM9ctdFmdmTbH+opoF+vlBeVZ5w/OIyFITEdmSAEN4HT/BQQFWR4lTLt
LIzgq4qedlYdv50eOOPVib7oMI0FPH1TsQ+cF/0usL2Xj01WXPAw4CasnlIOQbhW0miLQFvIZIUx
hHDRahj5bKVbh3rQuLXFCVfPZj6yeZ2zKvOAZZljpqYDktPqAQIXm0640QhhJuCw6QcrAMVAhPem
UrELevzIctgB7i9Gp/CwmVNCY7wV6wvdl3CIY9PTB319mOqFURCsw4J1Yt1uSfmrFai53UlNZP/w
mzYfV1Odh4+zmY4fUfrk/7j3Or3dpYVVYietY48WZEDE7LkSmgkvXKYgzBmi0+35GXuAFO08xWfF
YMO6dhDm+JrFQ7FptDjW68X2G3g2y2ob9YFg63CY8VwVJ7FUNO/piSNyrqwjtkDy+gx5oqMsA49W
33ZkLETEzY+9gBzMSLaZ935LIzWO1Kl+biS4fnMDhL4MjiD4Ran43hXYe6jjFbkUgzy6Zcc/n7UO
M9zLF8v28a96J+O9PaxIT7lOd5DyywnCW/8BW/7iyQbt9oiW5ZhAdIz1rw1lsmtpfqFr1nFwSjry
PJWcKCD/DGsFe5Cj7+ryWjW+IBky85JST+Vw81D1UIQ5dJdC5fFaXL0tg+iM2eGmxudCOFyg2QLP
zxzKnKMrei1eUvvMAcHk05N5bPbudVNGaVPjsmQDioQwJCpmq6DhHfsnh9TyJYFyCt99c13s4ppV
Et+kkLgTlTbJknQsyYwBT2AiEXn0KRAh+ZgjpxZwWbR/sHEyQ937uXHYPU2s/Ier2BZOnd04wkvH
V4QdeARvMnY6IkT4GDOBU/505OcuaihEUUotO3CwSY5Fk6899nPhJ066UdqPwGfilOXkmB0AdVn7
vwGRbCI1B91eh5dKeBZd+bUpkFqjeIYCEOzzBma/z+uYOO0kdAshdBjFUFNOKw/6QqEyX2xDUTIw
K26MdTKzgVKTEsJ4YtOSJiDrqEmN9tMSCjrjEKsi/7cMG75qTfRBCo3r0hKBI6Uuhci0tDEP0gNp
WlyR7s0Dle7gaia7X2gTwE7jzmoOqeoNM2u+kbrvVF1FYOvIUJA7D26+il8iN/2JOvkDzWn2KIUF
p9+6MsVuUshRkn2sJ38kCBPCtp3NVliLaDmdNE82qZoZgsEO1Ey7PTvjA7qCnMmMdknRkwAqmIcf
t73OPp9EPxhU8qPZ04Cz1vcNT8yUrR5bVF43lZIpT0iMjlG+yUUCuDMS/CpZJMcbclyDc+7jstd9
YMxe2oiGSGS6uWHryTxbgjMoAgfnm1fq2Z8VCEG0SRVM2QcrwZgMCmTQZWQN/B40ckIBK+yJynjQ
Co29ih705I2HhYi4PCOZ0taHWBCqrGclb0/tjgepCjTrPxOgzlJVRzeuYIT4VzPSu93LEydLE0Fq
TyhH2ekYDcXmTNvXwGykfPz1xwpS2xRcRDURrms2KqmMqAmWDRTrUNcUsBTWcQSQu5TGNCDo24ml
oZztPMNQYpcrkYE78UWR9Z0YpcUdkMptep3gcRnYTOjFsBrHbA0S2Ur7qAn549wuAPyUOiq3HjZP
3LBNKa64yBXbMTv5SqHtY++20ItFs/tS/Bob3OesBd1SUX+um9niZziJ5MAJwgEaF1Tg07ICLkKF
gfLsRBPNeBzVf8TVCxkf/XSyWLtglAelPHW9LwUzV3PzMr7GRmC+ODSelHgvsrSkrFxVpiRl5W51
Eqv2Io8W+W4OjcmHjqpKAefXutSs1UZ8ATnqI5Nd+c2npllKiUSsCZ4KXBo9p7CrvG2TN2uI2rqE
4HcBwHnpMVP12bS/lg8t4ZFpSkuCI8L2qi2CHPTlNufTCeYJ0DQ0oEJGINfeSTLFHJxpNeN0hVm4
o/AEN05mCSLYX3DidagahF2jPsiNxh9fsu/P60TgJYYbJaqYKHK4+nzc3jUAb5hHPmh0Rgkj1O7r
GhHEhKyQkjr67lamQxSHwDWU6hUwc4skqBBay5hp2x5anazzlxxQ+DDm0OxXo44dlyGpm1A1hm+Y
uoblyOy6YZFA808AjM5N/2DCLzKA2+hnt7AMyIOTRQBmn/zpqzqGIgZQfup7QrXyP8UqyjyK8afV
T3LPayPY7okoI9fGwlaMN5xYT/ffTnJvPbz0HsKI7c/n+9PGbzXiUfsVBPdfe6sK2y7JnNZagk/9
ZfpYdh7FNFFPWXme7WPIVBB/zkmngjDoq0AnPUBah4yq1pidN5DtznQjWUQyjDQQ0dHKenfMMxIR
NUWBxc7jLXtU6bX0JNPoe7qfaNuxVuqAqAy9ajcvV+TyR+VC0ybtDPkWZggbKvfiylBZ+BkAFeSd
0cwrL0zQgNvU626IN7ECNUCCYzcapmNYQqQBv6Wv0IvtPbrhjEn9NVi+SEr7zER3RBCm3iiYILch
9zKhpzvrmp2PaqktXbV9sOhSGuaXHt5cMywKAMG7dTBzfq00X6NRG1e7BpdxFuykZFaOcf1rfE73
MukTyiTYEgQH+tHQbCIoImcgiVVGdLYDBVExXdtDGBv+FUMiobYnci+EJqEj7kom7WVI7XOPvT7H
dbjrWZ3iS9OuHIqZDTgGlXdnuDQIbAZRPiZ4ALtGUXezPPOTeRWcCLP78sO/Dyvptt4hxmEe4BkO
6lyiOB8N+GwlaUBzFUm0lP84PwsjWUr2pezTD6dCwnvBmwLxBkEgeOd3C8jlP5PJLgCADCU62sJO
zb/+rZBnRPhCkIAKjOjguZ7fblH8cLD8ePSG62oEsjRATexG7WMmXOvUaf5nsPzJvMNKfp/MbeuA
GZVdWHTK0mpl5QOUDkHQ7KkBvxceUNgQsSP7HLs8UYHdakJRCxPPrvo+Qd2VPJx2SR4NgpvUsSrI
nBVh3t3TJbe+xP0HrDNKy8/VYTItyNrqZqvJ9ANnqAmVN1BYd1A0vjtIpnHBfsjkTzhHCXZy2RZx
3AqJrXI+2mnwhQ+eN/L2OHowEG5dTVqPx+PWK2gTazpdNJXNNJeExoK5YWVsbg4Dr/I0wqt2URI7
ekpzukIp5JVGbHxN8sXSfxw64XCxImHQt32uadCPHNdCnxIj+lyQrQmd7k2b28p2XFgkmKDxTov9
0oMZe4QP/KNuyNpUiQ7C39t6GDk4pJiE/dcwneQgVfazsLU7Nd7npFMfQM7823hTgY1KK6ASX8rb
Lv4CClUBYnLATZUg5g9uwKQGTarkde+VfjkGpDpkrgxTTXD5Y+7futSZk/qpkpEBpyEJ2QgVcl6b
r31aNZQOWdL+zSbANyi+HU36TosJdnZgPdb6OZcfgUCEVDrdljpeqa3QODRUWbZTYjXP5embUvrX
TMqj2JMirg3yEnmABYgcbBBdC0plcMi6VymNRu09zX8iLlGROU2fvUz+obp55FXnmPA6G5Ls8Ta0
dYuNODOkQj2OxM1xuoyXmij389oy+ntOulPwKHOARlrPgmW/WN1Qc/KL+Ce/pS8W8t8O52dGAFSt
ZmOqJDDC3JA8Z6sQo8wg4OPcZHAtuBZRaXcxt1fTyjB7s0yS78XG2Egm8hzz/BzII7jg41+Ii3DW
H2nQKWopOSJPy4azt6dMhtv1ZgrdrVbvd976VEbC71iFUva6cwc6kDPHWVVdXbFwqozCaZFZq650
tljEOc232B1NAR097mQcLmxbl3ALrc0jufUAeRuNRWzSD4ZF9oUui29skVQ+4o2WUqKwYIzMMCSC
4xx+Msq17fN7AvD++NRZzJV/LdQ39QDy3K5JyvDLnMciX2d2Q7IAW4vUUzjUoNVMm4bn0arFumcg
hgnS5l2GaBSRN2znYzffEbXUvpePV0HgjExeSSVdGDRAjb8SaF/FSqhoyyCIfJK+4gAkvShinHiM
U/AQ6PcMhQsUZzftbep74IVJLyaTOEHQzNikNv1k4KY6SHKy/0wOrZi6SrkYEV0SEL2QmEnSJWlk
wFwRdjvOeJzE6nM/A5WlpXZYYTgqQGZPY3JWAGSyRnjKfA25JeSQjV2/6hrvw2HaUcAuHSFbsQNQ
CSkZ+WEUW2ZgdQAUTK1UEQTgBhgLj7HK0XLuiac3Ie8f16RNUcVX4g7D7QQWZdz09yb5nx9qa2DR
u+bNt3klVWMQO27bA2dFgc7UUkHIB12iYxaS7rUtxIoTRE9znAkYJn/5J67+HD8KNWshtzUP40nY
dflkC4RnaLiJlQpryMNZxO942o+8oIIdVeGlMnboXX+1IzhK27/Q1Kv0M9RvCckjoKNGIblWi01c
DBUMervxkvWO/OqvVe0we3i6I0MCsOx4lawL8va4/CukljzxCxr/fak+Hj+asQsJzbFnn7aOgmGR
MFaL1AS2W9soV4oQHh3tQ2DA6rttoSF10ejyK7uLZw7KUpJuhq8DlLUQT39MVwwHifq/rU/QN3E9
zGUyGLdYYPLyFkQENBcmGKL1hYDVsc2C2riZqxbscTRyWLdXDwWRAv3jkEOR24SOmMQRp37CQJ+W
TgiNEWI6WHjvj7UcrHNLeQQuzX6xHmScueY4al4tXrtv7Kxe3BJYLlvvhtlEmDI0FA7WiHIoGWC4
NiQpuxfjHDPbLUzM7Owl/CSwRwm28fQkUgauk8v749bwkgxGps1ctkbgw1vyYyoBZh19GKemNNsE
k2f/ar3HjM1uxjIDokfP6o09x8zlfMb7B0Z3lMUz8LHUEgdeWH6AVk4RjKa8mlBSiPqUNBcoSp/c
9kWiTwb2cJgjvOHzCt7wWgAnWtInM6m52KmVD7yWx6n0wf+zmfSMhzMvftSuTtsUqxbymASDgRwE
9M0ad2gZhhLyDXi7BvPh/GKmce0DqWvbOpM3hlL1RzvXGCJgyYxg+qg7ViF5CfTqlNe72h9Djg+w
Q90/v92zFKuCF2jWKlJa4n07Hbf3S282cM/umt0AXY9FVto/gFilQ807a6cnwO2yg5uz0mTdKn/H
GrSkQ6Rdo4tk03Jf/PB6IPYAw9CIaa/Qh19e6drFpJWzDYlKgU/gr42nNkijZWleFler8D2lXyQa
4h1KXWViq08I78/Z3L460exTL0yKyiBcObhLWD2K95FbXfeam7fpw4H/1JfYeIqHgUKfmUlnayNF
EQquXb459idR4K7U7UAaMe+uyi59T/f8gdBTB592c7+65QFdZlgPsqQ+vnvK/2o1YQ4bBzsWnwn+
f5mkL+YXWhUlk2I2Gb07q+CjK+u/vLh1JVUtUvact3z9ihOYTQaMkC3KHAf3bxIp7ZwwGy1MkoLZ
EtHqLLY51J0BZnQWiigLx6m2Twmo9qxQrICuhz4A1dZd/RpVK7bu/2TSTPQZylsrsvIxudcmlbUv
mGXkEgVbXiYO0aW26RBcCBYx2TQnMevrRTz1ZaRtIK2YdHplh234jrgEMMYd82/MNp7mJ8OU3kTN
otgbTac17BI93fwz0etTqlgP3EK0jg7vb49QKt2b3C2+2+D8+nvVOB3DbG9doa2nhZtR4mILpQSK
myzHMNdSIsIuPa9dPN7UpyMR4PNWPIlDAL47E4agaSFm5/9PZ2qTa9h57TQ5erWCSU5hknUHjZuw
D/7GD3ArWTithuJZEmWgz3H3J0bm3/3rQd8Rclu9TMtcgdQw2/8eMTGRiA1QpNhKEj4GHGW9qQTF
W1q0jmaLgrN59Ef3hbDdtUv7oTzKpNE+K6RLpNwPyd1z7BnU/wGy1dVFlfHp3/K8a81WZjq7/w2T
tMP9q34ha4ySaGZUXajDsTbFtYwdwMztF/1EZFNd5j24xbmpW3yZKrJLLf8kzSNH6PA86RhtrJI4
S+1ALynirUBhx3oal8hfiTjzHe2GG3felMFlfy66C5hzBceoZlZZM27gkQV439+gE/dThQTXgnEs
cFsjzSJWmh5XQryvKSKr3USwgFIgOXD9OyOQm9kGGX9XmB6O7M0rppSSUKVvvZUzK/ME1kAl0XfH
Apqs1Y3vVNG6xiT8Mc24MYK7kl++yY2BbG2zIb1hzHKLyGF28XqV5b8kKqmDY1m/8mYmBS4GAXrm
QY2/Tl5gyZex66ogCCXi+9toCCoHfl4U7hiCgeP/78pFYnQ0SwWqw0BK0OOuPWIYW8ebwPWH+ChK
mZ4IXGjDsZovYkHKJEjmWHWzOceBBmEhmPNguMxziT2uwESX0QlllRcL0LxDKlx+dvLo5tHaWlig
1WgAc/cen9HtObGL6/TLufMHEEwjB/7il5O4B3j8iJ31KwBvDL8iLtEshxnFBk96y+oYbGYwFM9z
pxA+ZbnRRxqzXG8kHmPJjWJB4gcj8R0g2p5YLP0iz/DnZ01uss13+b5paFbug8bnlnjxNzUTsnuZ
UuNln1QT9TlZZy1vticV/EAO4jjiX1Ahb30jo7Jx25uvccWpUZ4H72dsG05/kYu85t3+nvLJzRVp
RFy4zm3ivRtn+ujusv42nmKyvpDq/9jRffWYsAJ0WRc6jCLzEEBTkXuO3l34tAwjB6WR+A+5cN/o
nJnJJm/8HvPvKgxrcru1p4t23fT+K5Omqgp/A4hycVO2crZ2UpZiqbAvftZV/RYPDKu2M/MgL8Vo
2xisyz2ccradiQhFn4prsbHQFxJNsxN3ys1uqzBuZtljPqpvKZJOJ4/iCEdwcAtxYaiVi5pGVd+E
0JFt9LfwpNicbC0e6n8/dqhqovh5BwHI9owFv7mBsMNdW8+DdDiLUkavE0gB8FHFo6gknhEPqFZV
Q+DmeatDQNuxN2CMZd6EAutZ9i6jewiT0X07Uupw10Vg/m0MMLTe0y3UGddy+HgQAOIzDz5rVk3b
1vL8/+ECVdCwtuKyvVyVyTsp6DzDrI9HG10l+dmuEV5z7JCUV/Vhx8I/mUVC+WPMqHzQ7P/79JGi
66TJpnsfaB7xMRsgYJUfX/bIuekx8xK4ypz1MleKGKziJJcuP/u+YXFxXAXstgoMP/38g2vtdtYt
EgNcQnNvj49fXtCCdwHHrd0y4+oxFRbD39vX5FBshkXRL4XAO3MdyMV696NBQ1UhZHghSY1ej54Z
LdlBiBuvVc9DaRSJCzAptc7ES4QCJu2il5+VRXHE5kaPqonHrkxCmHQBniRie2oRESYSL+14rTvH
2kOEgkeSiYbCOWEdyMMT3jZJiCrXQkJFgzL1Pz4jj3bSbETS5LVNwMO37L9IB9cJn3ORMbqhWdf3
rX60dfI5PHIXpSdPwBZPBOW2sQtBFyEJCD9HqG7V/M+4SqxEozY3l1DN4b+ARKeM1nMgLNG/TjkR
lzzA6ZN5fCA//M4q3eGbnnhQAciF35eJ7QrOJ7Ogz4ofRTHourku3viOZhdyNpHLVtuCEUIQ0JZk
a0xYCCO3E+MnclDt60F2dBZ98lBeO02p1VPh1+QwVcZnaqMwTIc/mHpboNn+jUYbqPkS0a/u/xkE
DF3q4d3KlFqczsF2uDnJajWplUHei4r9AGspxEe0dKIm+y5elW+MYM0UL8ZK6AUdlo6V1mMLiwmF
QFsNnuRC32ekDzMORu0t9WnrLRdBN6q1yV00Je3nOqUE12U5B6bssqkLLW8MkFSyO5g+4gWBRpoQ
DTlm9+dqL5HYNZx6Ik7RYr2+FXRzqkxLRj3/UDs4IuHKKCIxVx2fg9imWTlE9+C/9dcXsr15MERs
Hevp801KUlWGLKhVMdsX5HUaaMRcfGZ2D0LThx7AFohbbgqaNWYPgJ7FxKALFf0qWIpi4k+wauDz
J7E3Q8X0lUjROazhYe4yjg8kCUXVT4OePf/lVhCjcG7UywQvPDYvFr1QnVi7VrOcDx32svVwMFIh
3GIcq5X1F9Z8H80cr0CVz55TtZoaKsec/sFQibwE7MgnYRTSmNS6z93BK7jN5bMXnr+jO+VFU0KP
pnLX/Zd3f7ARUhv/u/mF/6z7DubN+r5tc00pwkCYuVbYChSRKm1aPhIdQs0fKtBmb0V5InmML0KT
dgMFN2hkNQ+RLgTKhl346zPASJq4MeIpfpWy6qa/SDq1duVS/k0NseoHRVPojYSpBxJxE5fraTmN
DMvd+ljn4VTAsPr0rPYjVBIwwYuw1BZsavURcSdQ5JqhjDDDuEi1T0AqrSYwQk/WXxllcdSnsGC3
ZFzaUggaXJMM8L4Us0k8Qv+CUMGKypIJV71x8he+QrOqYJvt3ZmOUXpcJ7YcwaxBAc8ot5FskoJO
haqdbl7VK8QcWqzHsNUIjH7uWIAAgOrRRfhwsmpeVFwQb2DH3swBwHI7CYHPasl5EMRfOZVir9hO
zrfN+IID6cUpAcNSiE1QyR9F82ZzAzPLmJLYFyPgIEEo6JwZ5PvogJJac0C7qw4PM7VSFxaEGzmJ
FF2dJIqHnD6UPCAebDVcnjrD2XJBMkokd8/Mc2gOlkjo3tvLQtFs9xfUaW7ZA17TXrKuhS1q524X
xEKAKPzqD9dtQzeIpedh92AaXlJ24zoUFum5wF4JnQWlMzwHz0M0KuJk1DInq6SfnnLm4a7zAZak
fDh//Q5Pm1TJqsGbXhLED/HCLqzXwkHO8Ep+z0NYRnrGCDHGNgWypGjv3/EEE6owWUjOmpcOjGwE
AaI2TSv2e8RwyQeRoXMZzaZs03EVcy2F81Q9etTgnw9kNocC4zx2TYvImDwFNAIvWqcdeERBi8aQ
JtyhGVYABMJ/thJ0HeJQS4bt9DhanpWGtPecRrhjtW5rxpFuTHg5OOKMEHUWxdkiOwJ5ZR/BWF9I
voTUrknOu+OdpALJSIKurtKVKp+kFybexJkTAzsJ4DAP4vSlPOY06qRZxn1MdGYIQhvFBxe9qGyr
ok3QQP/GsDkSir4xzTePe8ZoRYUR0k/XRquOTLYHBbsPSXXAFLuTmkXWx7+vkg3HXtizIDbVzhli
QNxjxEn/1aN40i1G2eAgZsrrOXUj464vsi1f5Vske6ZcwEsrB9h4CwDcGaMfejuCtqLsAcH6BbZb
FDSN8zwzIjZ8AP6Q5+yyrdeDRReyegIeMn2HZ9Vsa+ydpiFcVUHNcq024aoW6lWZ57ZeI2urNawc
LcbItBCe9l/jxNoz0SrLn9OOUWMz3ul/Sw4iKC1scoZGs4g7DePg+mmSbs2CtNtQloWu4DEFiEwL
y8f/Q6g4VujZetyiW8VcT+WRju4o0kzrD1gfVXs0CTyYX3R0nRU2oIsqdYoAaIY59xHYDymSI2DM
Mvwz4vSNWtS/zCzJkHIcponKHNKfrNEm6J7WYeLkN0THFVsvxX2f1zgg/Ug3EY8hDp9X0oxYIdl+
uFsMNJq/EjdDHzqNhnSY28XKGjuRgveHy6zdUKgDFriBdhgv2JQK4PMe+/pinWQtwPyjXPX4/5GK
cluJUny3zWewdmRfW9Xt4OFMct579hgyjGWfNU0RRN3c7QmmPYuhTVMIjbVi8shwc4Aw+AYAbKHY
NsLPFImjwevx6rD+b933NVs06Usv0qK3m0wmvrVIeMPyKwBtiPmpbZRYS8niuerX9pgkUgPCwGXT
xnKkR95lGY3oGptr21S7eE0DaPw0cwSEogulS+YkdzC6BlKJlqOYaj0TlUaUupNi1HgaEeVFS/c+
14FIdwGx7pKnpD0Nb57VQ6EFdog7f1wVOtLtkCCkaZj3ZP8yDiecXxjN/P6WkOC7rgKskU6fwePc
5YBaUc9xo3ZYqZnp4rIUGv8hEV7USJJZkcA0Z/rJin1UzvpFKrXsLf6ADsnLlMHjZ/ipji7nSz++
ZH4Og5Z8WAYMoQgzAGRBX+3i8ZltrRciKvFVbUzrvyG2Vhmuf69F5U8IIdINaMmjC+q90GH+TsPM
M7fB+A3XI9MEa3yUMk9jiAK06Uws5fVE42lGSnFQ2MBfY/wVEr1gRrgrpOOHCgQXMU2vzMBurTQc
QbDRjuKke6axg89oyOg5B+Tx+8uN87bDjr3zewWBO+77DXJVp6wOTM/UtF9i5IqHfugHO+755ORD
eJSJhrEef00tU2VT5fu5ieSarWs5ofYfOTtBJxnwM0AB8ASAdzarG2XIMdCL7lGTdDTimCEHJU9T
ZaQJvh+UMMj5o49qmng71EFM1jT9onwwVqYTjNEdmojxlKrXhYA6ZMG/kS27Kp6XnrFeTvkh8yfd
5M7AUy2uLN5lxvKMoa2AWlKt3R0B7g0xfYi1RaWQYMQBOvVZRa6XisR4rn9pqdTNezHIRKfmGLEE
0XBzdeX/qnOhJYJde+2nLppEBPmaM0XZyESnuJb9/JfkBO4xMyWCRBLppVzSyoorKvlmIxyQ2Im9
kULsL5fQ3qI9tbKu63p0FJh2GaMeGAnQd5dg9Ag18PSciGFN0EhsZg+nwfzmhcBzV9l43/RTyWvW
Bn/ZNnGO6virHMfD4Vk2QQSv7+QvpfZV6I6LKGm8TSQHFMeAbj+KKXC9eHuND3ZgaITzJyHeDCXs
hF1yfZRhmVyb9CAY7oPze7JW/WLd6DiUaVik1uJase/dY4uEL+ddo4yf86SPV8lhKm6aO7C8B/So
u/XsnlGE0D2FbNQXmL+8x28P3BLoQ47ecSS1BkRlohFqUmZDx4Erk2vKGjOlC3Kyf7vrWwBKCj+T
G5WZ03TTkt2N3hUQ+JlECgfzSLXTPAhOmbHJnY1JThuQxN/6O7cK7uQ0el+9DV5UTH2kebIQh9rK
KyXNLUgBcZAsMbBJOs4wQTLte6iGHSr0XO+CoVdS3MuSXVtMgQG+ETfyBbgP3X40pBS4u/D8iKgt
uukBblukSDPgOP/0npuVVqdE0BMsmOe6jxKwRoNnHFBUms/lqVMVjyizfvvg9ZeofxOqrt1+Xtnj
PWkW7JcAcO55I9D2RUkyi0+RU1yovLyPejIRGy4p8QnemuzGa+DuF85ABaOCJcIvn89Qq4Thv3k1
AIc03NoGZU6P3EbxOPU2McHJnpIiUDCh/4peq4dUJfpb8a/V/KAt27XuHoL85zZwN6AqtmM7Kqzh
Y+XJvctNY7y43kVN/QIveBfkrppPA02gT5pS2FH5R6C1cYv2WyzyZl+IZ2+4mb4kXL8sVgsfxxuo
nare3Hw98kHaS2LQ67kimF2wJjsGTzV97LZUUSjvnBaP327Vp6azbF/aIyIfI1H1osmkhZsFL95F
zIb4EfnxZbYwN6hL5lLgAWZuDTsgxFUD+TLytnvhKX8SjrGDld9OHzxVy/Jv8ly9vkifqNnu7zFv
8KDbyvDNI3N3SISF2Ru34X+jD+O4zqWf9IxJJf/jcZpJgAd1qUwa6aZzGnXkz9lMKmwzGvJ386b1
hsT7q0/poMaIDw1HHnj4fRjw4knkW/SoZGP64oMlESeCegyC4I3mXxifLqbRGRRHzr1j4zhc7rQD
B5Hy0csa2zf9ZnHpOM5qz6medt67yhuSdC3Wd7VVf9o/p3Gpc9t7FkXJJxAESvtoio3a5YsgERf6
/oLAqrw4Q9CO+4u/ZohgAnUQkeLKHv6Sqzp+MWrgXaMkQCoXV6NDANE6d8jx2mOo2jiZOq1f4pDw
SibvTnUP7wpZY5X++8Ijw28PbUc+7plXYvIzsmtiqk3M3girtAFcxTxnDYLh9PNfosnUgsAO2kKC
3KZlMy4+4Vk5AwH5y5xd1wWVGcyxBWBuT4DP7+Wfod+O6bmpGI1GjXW1WUzxD3uhma9QlMGM78Ir
FEsBJjYoA9fNJdkunaXCM7CmYzRbEd5mrLmQ1lfxOY6tXteINxgt1mvOZXaN5T5k9+Ft+Sx2+UYR
em07QTkDD2QbWscK1ntQoJADGM1iU+x86K1+Zuw3c6WWdUVMw0/lsmhgNnSnUVrAMgBmmtA3i9i+
4K5Nv7OcxKCgYBfH1B16IflwSnR6I3G+eKJ23JrrJ2Pr0cMwFo8VV74pejozxm8kvTuKLNTJbPJn
ojjZ4AfJP3N3Q7KvGSan5ZT5+y+nJ4W+Gkkq3ZWed9KirzvfMxqCrVbkNHV5SxRzedUH20nNh83m
2ujOs070hD9VEvR+b41bDoGVB3jD5PwfGh+UOV7+p3MEtZVnfw4XSp7b7CEL+vPkuYSQjEp1CLHc
0/EadjbjBdLRzkicicKfw8HDZ/W7zm5y4s+HKLpWhBZBZm4jebcBP58iIiIBr7M5cfoxwLAtxA5+
qOQD67GLPz/qjIrFBes2nDyxLVtOHFqZdNah/m7RrrYNPrL2PvPDsGst60ExZQfsXAPUJKWdooWn
ZEoQCjYbD+kYVAj/UfxdXM9MF5n9AO5NgCeurehHLXAT57ts93psSEJvW05co/kusa1dy6ud8b31
k4iwK14Y/dmUdlRBw4MF9fzjU5CirP0lq91kvdE50P9zvULhUdgYieHpW7j1b79JsTK16YUyo4Wk
We46gnxUlwsFp3I74ew1uHhm7XjGTH3OeFkRm9rPOLXBubkyruu2ruOT+Sug5gY20bNGFNRTTULh
+zypBswhlKPUUq4CVYIQRXCql0kmEzl7Fji1mvh2pUE4SDHItp7JP3xnHSfNdyK0F4+YRQWTqFmQ
FDXFyzJhnKQA2qEstRetCD4RtRaHGcNG5zKtEdgOmyog4I1Q9GLpgWKMs+yLekFc9BC1YssQj0P5
rVK6cP7ncyoljoyY4etuW7LUXXpMjw+2MMlVXT+pwPP0Idio1d0SNXUsvXETnxk55L/tarOj2Kuz
E9Xn4x010fTiELu8iqv0rYzuj54jTEivhPIcAd9ohT/nv5hmEqJN7aTDI/LnwCEmFKkzq9hNxzt2
CNNo+REoTuQTqyfSoNLXQoR6B4lCbTDPQ9YG2jKJ382QfZjtwMEIVAUzE3ByVpr6AeOPWFKMB8cf
P8ZfJsqu0yCr4H1Pr8uwMZr0zpVy35kx+2lXi0sGWddESwU1fh681IY3mecVrBYyFcjPvsufZ8bz
Uq3nueBzj2v6JLs/a89mlVV9mG7du1SjI3fRfOWaCMe5RnXKPQ17ZkF2xXe4roNWHdQz6DqKjH8N
qzG2RjjNLp20GQjehKHm4Lcq34IT3EHd62XysWoOM/Y5B1nIqERF+lX+reEMIAWKIx4pOnpWsuRO
+J0/XuCufLp6bH2z4sam5+AuwxxgXSBL5slya2lckB1uFGWmEp++UJamP/OFEumU30UWy+rlq9h4
/aKERgVgReacU7GqmxayktZyBMkqfOCjSOzagI7ceO4c6zM7EJZortuTCg3tMY5Hz8PH33JLnX4b
9snShtBnb4sTSy0jMFvkBAGTNsC5AetALcKkl9+ZP5fBbHt4j7soYvESGqL2VNVV3bxUe/4OADLq
ij/zuvk2s3QSJqpxyJtZ4AZQGvnJcRkTs1aWINq6aVqrR584GZD/lBou1RnfVXRvxBRSk3azi8rF
ZYCwuYCtOLsyH3tzSxBqJAE9vWoUwNmmWju3IYQQzHPIn30AUE4OWyqpOT+LstbWYLxNuGzFx4pj
f+buuMZpkPhbOW8IE5NLGTNgV8DJp4zuEQoymCp+JTjLjJRp9TjPL2ocmXKNbL0F19YiRWTXYq7T
iAaKpemeL53gFVRQjCp57st9nUvqaVyyUmt/1YDQWMmoMy4f5eysI846azjd+NSOBI/a43tcYXnx
liUSvwfIJ2IHwq8G2jl7XSk5prL1f/l1sKMoaM7UCmsKYi1mjMu1eWDWmt7zioufvtZk350bW+DT
Vq1D6LQN1ZyIzXexl/Tr2GiP7uW1zVx36RB+y4EaoJ7vKNejmIhhtDCZ1dMHqQ+tn6bFCgpgJf6B
mKhHu/cuKoPXTsdqDYAKCxVlb4C9dtmeJAtRzZPIuALDrZpJdZOex0MKc0+YYChqz/zpgMQ2SfRe
tX8UZgE2iCkRSjNAtXGYHDvEaPUycmn7izCIfHS57iS4sVUx0t56q73IbNf+ek5cjfSLRHkfkk1K
twYM6juN/x/unxV3+ilHvPxP81WEH5b1ECC/8xTpll796hjmr0eBcFXTCBiKNR6k+N77GJDjK5GG
Lr0/pHzhP+LTa+uIEGvNeno6Uy3ykbaU7UJ/eluW9OVnm1cmsvjv5YfWlYS8cOuDjZLdynRYYMIs
+7PJnMoseZCFBBos+H7+m64TMeKcX3eG7fAwUQcizavHv3McI9ZU0UJ3uC07O0PVn1gi2MYrEpPB
o1ZzVcZjYo+C/AcbFf8VTxrbZ2ID8zt1ssmeUfsmhrHRSWlcJGStXB5BXe6+ej52kGGbrkBJ6EFh
ZzX6uYGAovYl1UK0x1Yj2XFGM8TJLeWF+ELdEkJBJWAOaBgDm4GFJtAUzt+Qjd9HHaF9nm0M50TN
3FgwL/pAwoJsS7orWhKlRSEbdA4eC58civaqGJUouW/jExFrSco4/xrehawgpOD6HGWrK5vT/rmF
0xhuGMem2Jj2uPsdFealrYtIoS8PcD79Ub7bJqkLgqK7+ewLKy1mF/NXHGs0MofhrIvD1C/0muv/
PY2R0yMuSSkRVnMDpLVtkcbTRxSTV5quSEONRjJczaHj0SWfMMQ7gdUPNopJH3WE+zs4d13DnFFI
TVDj+gTbGjCEWHBd514EXhKkZTb+nMof1iT44yi/d54oMBJR5rW2bz7I9Qba9Vuhx6LBWdc8gvxd
hv0z1A+dxjT6c2ai81DRdpvmQVUBn/kbpE90G4wicM7BGxlsFB0Rw5C/abYDLBcNtU25LzP3rVZ+
map8dIODeWRjL/UvUfKvT+h8L3uLSIGysr+Qgz1rLik72wzHY6NicnR7xEJttUMDCQh0tuEq9Wde
dE+W1pBRDsehTj5elQMRtyrNnfYjJedvcWtLWaQrVHiw+3JvWRnv3YM+k2vzSVMBvhCrq4HOT9WV
As2tWVmAbd7wldDSWDWtFMWZK+vZIdQI+ppH1J+y4t9Jg4sD8hxsJxwzUtiEyUZLCzgPdvtlgW5z
G871RErskLwpZRrhI6E2C6lWTCPRk/cRAEW1QrDYfpO8xalWlU5CD8a/ygRI5rfTycYjEgFp99ko
cWDSoU8P2LeUEfaYhjLtBIko4yQhx4olPXQC04OLg6tD3/kLY7ZLz9arKpEkDSQ3MU/fqeB8pyRn
v7dmMvsUOU7/1hE6bENOQN64t+tY3Oaf/yy3g3Emp2s2HOD1XJNwzF7lI3lj/xr4vvScCrWefWRO
9m9K/yRAHiB7ZZL4Xfq2C8hu9PqLqIqTq627SQeBqxf0fRpBGRokzyteJHknrED0r/CmAYnEV90m
m/YZ4GbY0WAtu0gG4nhUT0ObMyJA1bQ1Bfx+ITS/hZ3AmgrsHnx4qSSJaGznQ6ZcAJW16hvwqTX4
sRWnPYRvmOI2ZL+crSDEKD09nJPRQhN7iJ8jYofHOZtryCvZdi/xtgHflNk60xZjxyBFi3ivShsl
pAVlbmMxaYslioUljhEBnHaIYce5u/la0B1dxzt9YSB1CbJc8Q/wfPIVT3GfG4Uy5orpASu25c7I
P/TRrjunkKaZPNvbvfn6JdMVqAX47ZXovJyxgUso+7hVZRu12p4KPMcf29n639TjWhpmxP3ZvU2p
sIYofGwtnPsaG+HKT0boRv1ec7jM07PJpx6maMoPVS9FarDjhYq4XRKYU8DP5q9idre4Uit/44se
l6PdP8IsoWHxdt5x7ZNsU24xRKOGCMuZiX2V8iBT6AsTXxWex9ihoH/kvNEBOZUGnBdqN4dH36o/
ieRa1YUBfUUy+2G4qx4jUNgibS/b0ELbNjUwXEv085Ellu8m9QJ1P7ACcdDFReTkw6crYHrMCMRL
oX0ff7BbmH3bB1dPEhYMBWWzgbjqdwXyx3SIiBwXErLU4se0zBQcqwDLlWgFUkxvMb3h7qYMusFj
DBxmPiQEAdI7P821T0wM4OvN1mUlF2YjrMT7gv+aFREiCMs4qSyLT3viMi1qljLxBd2yeVaagtYb
kwgKh/0a2J9g4/yGrAtSs7S15xAJk7btu9x8ehEIn8ON9UIyDTuMDkKtk0rsoSPQ8vZHq+eXWAuQ
BzN/XByadb0C5ltw5IEjhP5T4FkMwmfRXd0rwKHwtf+USTNSAplW9ZwOKebaFH2iZccQUlTe2cgL
ocseYjCI71rdYov4LaE41DZNr4lnv3fyrFoQxA+FOQ5caKsdrH7YdlC2jSLB9P3HRnNJnTcBLBV4
bJIND6NJ0R07Xe4d6kWdgKy3AL282OLXzojI2noWzbRIgNczE/PyZNLYDShORPo4V5lcoM+H3LhT
FMCK7sg4d2ZNO8Cs4fBqMNfOs+mDPbwESfDEy7o5pC+fDQTH6XZrOo5hYkXDSkPlPcX7IiiycX9v
l2DqVd/7cP4xKPPlsyZ/eJqKpGhgzAeZiCtS1RLZHwLqNooNqhvY9aU/Jv60mt5XP2O7ZDqWtG31
gD3ykA9WIQCNqopLh8E6q4KC3Fs3jSmdn76jHgn61Eqe6qLdr6IQqSXD7G40jKLytuoCF4sm1fac
9Df/UKFgRgFAftRfW/xNmZU0IjlJMOyoYPVLa+raWXjYpCHih04KoU+tR1Mv6OPpuPytWNqHucSG
h4wcbxHPvtyPdR8XQ8Tp14qinOwOHpv/LlnKPtznxScR8GLMvw89sShMzwEBK3z0/s/W45j/9f6G
02XC/iFQD873pu2DPyEzmy2mUawO8aNN6fyNLYLXHkMFWUd9aedbhDuX3FEyk6SM8Az2rXH1zJnA
51VPGyIzUt8XqAJ3ra2yJ7v9czWTGRKrUx5g9YX19F0gDrvc9XNNot0xvCz9SVdgvYsK+dCpH4G6
k9erAWWfgF0IRBifuZDni5co7kxQhxp5nekTe2+yPmJex98ngeCPjl9J0fywZYTh4YjuMY8JsQnn
pRsphExzl1VJC3ONFcR0Cja1PFwBMqaAPfCtAGI+iDMBrw8YOeH8j/jgVlSqojsZEFIAg/r2y7RT
c/vZCXBe+oQFPptPHG+e0QY/MXKDTQgEp/6p6Ek2ZGq4qXfVbYJejn48kklhNpK5JHXk0hP6BDxu
6mywU7iTuhP8vA90Xmr0NqLQk3sSoPH57JcfST8ZuJ5YK1VFks0xxP+fhLOxVj26RHPnJkxScu/d
2KEZG/sw7Crr1IllR65xVIaFntge9FrfJmGTqtii6lJYVG/UAz+xlATU/yZgd26ezZP9QdHlCxc3
ZqV6AAvXvhj3cLminXKJggvWmKr9iDKy5mlZh9LZMlNDm5LiiWPKEXe31A/HyWaIVKWxEhqNyHyA
GtSScppiEakU/lcRTlxzZ4t7405uo5Sf1yCGcMo9hgZKiZmSdQj4jWytmvAg7/fGcNh72fJW5MSD
lBOr5w9g15z2dUsPxcdCC1hh+TV4p2AkDvSZ7jdRhZmD+VUfM7l1TJpCrcM/YtATra75gcbaGl7o
k+OLoi461A4EUTWYx00YcYdPpdkiWIxQ3YqT2TjkMai760VWVLCpnhsK46OCm9HVcheI0NbUc3TB
LFSGu/QARoYIYuKGezhsjYW5U4UeuCysg08egQOu5DgHhWrM+01D5RbISY1kmtJbQ/FzBBsGbxWa
5wzp1Qm3UvzKXoihqBw3yA1tJL/6CMV2QJ1tswqA8aNVSKB1XeiwRzsfRUZovzVribco+zoLD6if
zU0LvzCgTc0jNRQVZwhMRV8w4i5K5Qi9RdJwANSParmsBv2rijSi777bB36GrjlGy8oVOf6jD0GW
e4g+PZ1cfFI6WET5D0pdyoFeQ4T3aKmMEP4Dc736neYIT5PeAZpjoCGBN070A4Fz0MveNHPuOwXP
4P3+hThwPCJreGyk9PciMrHNYwQaiYk6+UFLRtNMyjlqIn6OXvj4xY+w7secwgt7iBB3WRNmA3QI
wGNZh3+OHKyx9aEWCjdAn8XMjXargt1XQYOfDNNZTVBf0tl1oFERCMB5mgxpZ/OCt05nfhOhmUa2
xgyhVcgKk5tsd6fNw3R8YpDtywfdKKT4MsPasgJaHX1l8zchlWjWvpj5T+XEpX39CL7sY8DS83e8
JjV4tGT2tMSPfo73BqL/MeC6uPq9ulGh3SMdoD1mJkK/aAxlsd316/UZ6UUNy+bM1R8LgwksRwZx
zZA9561cjdefHNKvhh0bNIn0Ky1dX77amgNwDNcHksMpqSYkkryyhw2e2ebNFUwYqGpGUZuYp8HQ
pO/MbgfaTpsUDcngm3N91lTQPsO4mFyaImL8er/IsNkKJA3hIS3HpN2AYlQ+qx2dI0L5Gx0pyPU0
Z1iYs/ezH9MyBLQIvqwgVM3ULYy5lWtIh7I4JUQ7x4+Iu6+fIZR/2Ms2wBrYAS1R/JrcvNyElgFc
Gd4jUfrxEpWUUNjl/wF9LJj7zYKSf6kBNQCPRhbcJNepCk0fmdd5dyTG1t5apbcbzFZ04hygCtbA
mmFiARhek9/O+1f7s5DeBzbkWw31DpyCRl2dYJYORj+9UtP+UOWunUlTEwd/UE7/7j4gKN3G9TUV
gpAlIjoKb9SsixGOfrIs1WkznsF/W3/bFA86B3b9YFtpvA26JHnU+J6lOJkRvZ0q1db509xszF7v
tgPhaaBtjT8+qUPtnMmydlWnRD049O6xv2V2MCjlS2k0lqostysDREpjkoPzgbyzqXCV6xJ90upS
4MNR0gmXyWJ3ov/2LnLDjRvIujzBLNYr7qdYAN14si4/KRExn8qIdilLkLkeOxxZD09RxGIbaCs6
yvWAlOzCOJ2/4UMkWTuUuEtqxYIhZrJVM9poXh9VTf4H0OJPGudcTgMAwpAeVnsRVDKcijpp8Kb9
TNqorgj7MV9iM7zgIlfwU1gqr4X/C/UvFzPEDCRo5RnVlE18RMYvDBcaeun0fKaAfI6kwRiBPi8B
9uj1Ihc/FCjjiZcjs9mxciOo1NEaRI39FUBEOvUIKShaYwkVzRRQCSnWrsz3em0J9oTCIjiUHzVA
K/9KZuttgSBlwRlFsU/6P9n6xEwfHee8VDzvNbZLdh2+16VYBQ83PbhcbU8zjnlqfCieCzsI3GwD
VP/LKHAHN5cxXBcf7ye2Z6BSTomYvbGVr+e6WH3/ClxLTq7yw+l0IuGhbtyBczjT7W1jbFS+z1ln
FnlvFoCgmqshwiMolbg3ylML/Djhe8orIIUHj6Cu1Fv64zeYnHPvr+2jZaO7GZKK9tn8LBidtaFi
EHMa8ATOME0Z1PFVPLfjYTiU6ccfojC5OaFjlcYn96QjoMDZfT6Jk5Dfg/hnQDXtY4Duet0caFGu
I8vK58c/xQqQWr/4V2VxK7dZ9wTFsjkir5DtASIKk3JRKW6OS3uE3U6ZTS9A/ejuNYepb9o/tetp
pyU3jBDf08U5+/dF0wmIHbLkhcQVlveZtIqVdmHidt7d5rg2UuHoNwczJZazGtNUKnEoM7PQl1Z0
NP7DzKo80p7za1AhtlkMzwwkFcJ0vIgoMh3rwKkJsdHZNDfUw8MR9nalW+hjIxS+RNUfvJbzxKZT
50CXRhu49elBk9TuBsqZ5KOygRHRf5O+WbzkvRnLB7ou0vMSBYa8IfZWOBVTbrL6jmvM8WoPsJ0f
ayVwwFDB9sZXMi01THIaKpHZ7yUiAMd9M78fuU/g6nKjblTcg1Pf+OVCbFIAP3QYNNccpUw2hQTR
OwFCRpnC9jcxapL7bI+nVRiP3EHWBaBf9PmW3rwLSe/yEIfXjA0cmOlYevNLmaKSPmEjC550ZtOv
7dMVxn26cjaOK3kTICK5YxXYD0bFZFAyuov+1aR3PnqqFoOG4s/+JeEIO1vrSiyEbR+W4q0kdJKU
icxBL/XBy6ZwLZPlZW59B6OPbm2Yt6KsMnhayt33VA4Fy7myGV5SvsWa0OSa1TYlrskODwkRR8UT
3mNRsQSZZ4K4tbf0k0KbkZ6/vptjupfgurOSddoy5Et3UWoVjdStfr/9AIbg0SAJn+JEswH8wi6G
eJuJtmysGNIxK3PkgIEsbiH2BbYiiT3YjNBzjqBPPsAeybWud4IA3Kj8RAQRe4dIZoqQKhrZ/rcH
j9Jf+gLHTTnm+AG9v32LlHFkla6w0Py9QYZDaL/hOd//K2wK13/MKj0t50Bpiw5Sf7UhQ6sweRmR
fhZIjnXqHVTXmBfUmPFuRnuvsBwg0iSxrHc5Mxm0Bh2iq4aMdzYZNSRJ4D3PcQyZfOYzClrLQ5pz
kFdu7JVAaHA8StE2fom0UNekdDfiwmkAqeDvYJ+jMI8stH7fN9fi+CurXtixbA9ooHx+8k8S5IO5
/zALWOOMGIzxiJQvWaGMmA9Z6raZEUf6mp5koPcGCDqPaoVmZ4+5vfvTDyDTLpArzGEwvxaTfDo5
VJQn9wM1MQeHuNJVl9doaq68cYuRvs3DzNbcB0Nv2oM7FrYerZ4PxlExS6uNh8u1F7zzxcu/afEX
p0czR7Uyexg9CDn0KCALYyonGJqbGbvw3OZlq8BPa5fz/8GPixV0NOQxRgym/Ypj1dQwe0WmAFvZ
kkRAsGVd4c9sYIAwcFcfNyd6K6aja1a2rY5+yngrguFyq4mcbwRWkhrY7KCk0qQWX9d/IcPClyoi
XMGwv5ThHQvGHJWeTC/+KppF3DnjHFic6p4Ka5FhPrJ7OVSQgOJ14iWYJ/niUUf34fCFPb7Mf5t8
r84t1k5HY2A3B6wyDAoSis43zDLQ6qHp0g8W8Oi6NPl/kLmwECAPTR8JuNKIgWLB+7gUQ4h3+DiW
Xm2LbMRfTPwX4bD4RVug2KVEeuXm/hvOFLaLiHhwq9frvukZ+4WDytox34Zd5VWIVE72IvSOkNsL
eFHRfi6UGIdjn9/cbUXmWMZ/ZFVbxNjzXYIKVbw01Tm25Dwlad5xxZqDX1T7hVPRFhnV0jIkPmSH
DCkFxwFDPTJVNzcEhZr/GxXtRYE3idcKpA/7Jc+mhHG1zKo2SWn6BTNzd4f0gmK6tRT6ae7B3pZZ
nEui8xij7TW+3dS0JQsxdOC8BmxkLsTGsaeVKDDPL8zVfivMhNh/+aUXEOUVkHHHXeUQq3vFJ8s+
0apzRzRbNjugjsak2/BJf61WiArr3xHx4NjAzyQoiDCBgCo3Si8VPjTgjiDFWg6BuFJdXQjmUHqk
ZT6UqzbECDN4GZbBKlF805XxnYDXb81//edxHZaNelpaJjWG7Q+f5msRc5fhgOr3QJ5/lY2kdoLT
52QTCSumOUAQllGisrQc3Ok063lgf9Do2/a9IScOwKOgKz7t4ir2t6Xf82vaMkP6DVReuxHNMPDN
LjteJlgNBF+lDopp7KLgn3b7d2/DkHnwL17nSfGPuLh2MqlZpmyyc4uHKEX9VRgbHKE1TiQ8xGFx
LpOfVT9AjHpVoTV6Ff+RpQ56E8WeEawV9U3svL/iX1P06HwItPCm5tj4LH4LHC0PqQJQ9ZI+MFSV
o852WmkMPphtxnb+DvXAGUEzOeZIomSp8sZDNLdc++M6UGldSk1fG8LTMx+hB2bEATV0G9Ll2A3y
r7pEjHRPW9f7gg88+NwlYXQsKKXzYehALQqPpDIMQpUOG+eLO0FNT3p3SicnCYP4insSi1zhFEnU
aHj3jnRNtHL9S1B4BY81g01u2AHmA5uKTNRIzTEf1xXcZPsoXVZscNC7qXccDQLFr2FvyNsZkbzQ
WuzUX98HN6ypuqT+pM3O0cJz/kquz7mdeLAzgBvlYAaKfMAxkFS4PT0EfCZKJFchpHl1Od02XCMk
XrpHsRDyQoeplBVOIl/+yN2b08DyYWGEY+4+CsbxDEboMBykl/NIweub+pm/4y7l81KCkFtsUqsZ
svQkC3KBtvne4d/dbw9ooaodTedG+zrPOG1BBcdxvHPXjHi87VesKhHgBNReR4X/UuLKprwtC706
lMRTQb+3SAASy/+L5+27NkuLMufQbPXX1vMGWhl9gniXcxDcYD7a/FfzQzpOSxNGVWHC1cgr9V/0
/Erk6FU9Ow9XpIt01fitwR/zLewKqc4DTo7btiS59gjUyyjELY8K5Mj1b0ZfemKt3QlVaEbbOa/0
MaI+6iOq3Libs4S92yuxa0QYPVt5qq+Cd+AvgIu3ATROFra1iMJlTVYwmMcM7jUrkr4aTbm5Nroy
QFIsx/SLCDtkg1dOeh28ycBvp0EMdcdrhbCKCXEwg1ih0QQWprEX8FWdTCOCRXrdtS+a5iv9PihV
pmZbcTmjAF/+eOm2t4siamFDttbYd97SM/wOJssYpZBmiH/f8yQuHbfAej8K6bDMQm9NG8pCICh8
ZUDI8o75aoPKqBEeAVOTv3fldosLvVN0LCynNEzOkI2jmP4/8CWpjB1r/3DnCDgjn8AQpgqa1Gfy
WJNsnG5hp+bLVskcPuRXcoA3nyMc1mjjLcRAwsbw65vZwGM+jBfu1KudTEa1V54pnTBMI298YG1A
aa2/h0E32j6ntwDb/HllBuXOF7bwiAP5xDsaPpOFgylgDhP7WYJRmizhrTm3/2TDFooia9p998wy
mZzr5kkHXh33k/tDJNeMisff/Wh/kKrAGq1YNUee2CAu5zlJUgjgFP0Gp77LpUGmIPQ6imPg5XLK
wn3lhBMpuOCtAzGA1AN+eROoPLeoEYl8inPYDo3bGoslKAtiFDqBUqIDLiyY+Gv24DERGYwSLoBq
pTJdGdccju9OaaRJtQ58YpENwJl4edCS+i6jkzbrw+oYDa/LvDPLiCEoqmbF6BA7Y470VFG6gkxS
5ZWDBh0jtLd0SAdzdxViQxJF1y/szAWyOv3Ja6nOQc25PAO+ZBm1UnV3rSH+gAyiiIWvCreR4Z5n
GWvAWIF/cKNNN22q7qY3Gz5fFLh5WKS0RqtJFgJcPtx3eNbZq5ylMl0T7l1mYhd7fZ14WUNHv2LL
Vlp6aiPEEvqGAF0uxBVSCxTmgbKJhqqb81fSFKS4yvDK/l4JFoEJCFsAhjb3+LmUtT6ELGx395hE
iCNTrLT3Qc98JED7yJxwxZ62j/fhf0LR69UyKBIhi1ufACKAd1Fw7evt42X3jp6n7G1gx/089zl3
+MsXLJNRzyK4y/+aocqTgZj9ph+UENliV2W1MPMFeQQLA7H8WhOjbnkkLRUNX4/NUWBXrms/1z4h
etL/UbuK6M1NZvteeXgs6Swx9h29SJaNquHJ0NR2UN3BzPbFtRP0wGrSFk5GnEURPIRJxniarIcJ
sDGqZ3WeaRh5HFNgysAqMwN5nrEtYjqFQDbn3HKqw65oOIIjLObBfFvt3wCEjpNxqYBcdMobcw/L
lKrK/jLx2jOl5d8d3QGiylMQENParEc2AioUvGiFyoc0UWrUhgTucikwor7o97QL5gHf9buD5XnF
ZbwX8GsXDWx18yT48P/yu1aAcTZdVtBaqiQnP5O2dbIFE7itOEUOYn8SiSO82HBKXyJSK+zJfmkP
H54l9Vt9IwK6PuHsjnM5Ia6jFgbzJDRAhe+yBdOBdrUHxZTjVCnPFo81Yk3GSLKASmGb21Y5Pm4X
LksjYcPqdbWOnf1oELhttmFp+gyiZroXIVMccwP3biQZ6NddN1J7t53YNFlxQ2b5rvz3PY6PyX1t
/Cvpb2kLOEZ7g/qwUrxCvqV7uTpeTSQpJ7uj1NlgnjtT7gC85wCC/fnUp7VwB2XN0vnmQtk/Zt6+
VoZN7mwiyNwrdJy1fF1r4XL02L816rTRuA4wkgP56zjWusF5uYw1YKj2UR+1Q3sat2MoF3Pkv+vY
DwmYnbMhIDrPwMWJ/SnsYLD7lTm7s/qC4KiPSX7JBgF7dh6w1GKB06q4BF/581pE5nuP+pSBVAth
h4lMtUlrcaTo5p1kABc5KkwfE3X8YKLzBhb6pYHMv/Sddy898P5bdaKHT5hF0/W59X2WokuFZXu1
lBoLx07Z6L2u69bDMqS97bhQULrf65YjbyqMM1Gj07tqIhM/JAnRr1iMVKQzn/gPLHp1He8dxk1x
cIL8dCyTkZ0GMwk42Gwtz8E7mTkbe2SDkiUD+ebSkw4oQqN9qh/KcrA0BzCq9mHUYnsggC9PkB1A
isdkDWNWBZejwhak9FHX1tnk9BLTxQAhLPf6vnJSTxncppkhLe2m3r4o5Ri6FfYEqaV60yohZaiM
TTibsaw2BR5ZGSTW1CqeNGMUN+hWP8zmiC72PFvpUQbtYTDKvVgoUPdabztTX9KXe/dVzg/2W2Bw
VKr74pLEgovdSk8lS7R8cLaAz9R5smR3AAZDey/GTDV+P5r0qTfcla4DkxBS9IVyni/qOJPhVCep
SZNNxG01kUNLQkvhYgoHFrpLwKoa3cg/YKL59H/1elobbEPTPLO++5lDfr8HZsw6xuY1lPOJbTux
baZV0nDwA7j579KsFMmgJsGb75v2mdMyrpImlKkQo/Emp8P3kRflJFRoCPEeT3/Ksp323tXDKSLd
EzfQYJT2fMvQMCB8LwNvzW+432UhktYpaa24iHAWUBu5fzvybjvE4qQDFx8AMuJJZknemBLy/+ku
qcq1liKHd9atS9ZdLnV0Q/2NmTBcTIbwM6TVhFD/lDO8VJ3EpP1LbteiLNMHduy2hHlTSpXOMit6
K8juhqJqG8eTDmxLyE0DB2t+xgMkKLfWj2DrI9w1R+HWk7Qsyv7xKE7Nus2MVjyEf1Y3aWW+04ZV
+5geSQhGBEBV4Z2m00IBW9/DR2hkLRG+Wx19EhW9WP99P27zHXNZbK3CdMY6oGQA4+/P+5OvPofR
IAxBJKJ2QNzKayeu/6nHGcrUVzeHXbeY4HoOdRmotWQFgM38eUZou2Ic2J9YO0CP3opjYDNzhcfU
rv6c2wYdWGOPQqCd+sNwZL/6/YZ8pxAewaic+s5WYy7eVn5Tqq8bPGd3Hy1ReK0AfIvVJO+8BT9D
vLxHG1VZVtxaKmf5zfcWXo4HeI/+qSAvRwVj2cizrFApiZIgjGD7s2znFl9tMhbq0aCfcXjOweDc
waBeIoNnmWOBvsVwqJsctozzci3Vw3ON4cNFficxeT+pqCXnXEFe6YPg6PxTwYNq9UrYQjI44mcf
1ls8PLPBviSWw/SlwjwP4foqoy37kG0p7MSRPYn3Pp83owDtHrBooquAoVxSjgFyfrLt10r/LFcV
/TJajGULrkWWE5TviKrbjlD6AGnMp1ydqD+2APappaRgQJSH6BDfiE0hoWY2svdryMw8xzybw0LI
D10bKLALNtvkbxe3oUUK8QJCIH3nvk+tKTqDlwigsoOGc2GME+AQ2u3evy/fgD9VSnum1/9XmbHK
XYZUs7cHphvh/lpHvAJt6OB+qUqd0qkR69fBOOzOLuyx3dP92tC7d2IBwz9rZ+/RFPk3Hl5JgfVk
/qQ2NxwbvvX4hfYoYe7ZWElvQX40dfLVsM5r8ylTuePEou05qxJKq2Ytktxlnr7djLzS/ELih5RD
EWMFWuy1hDjxCameeQkkrF1CwGJVxBnXVPFszUrBiXH1DF9OqUGgHhNdmQ1QvBVdK5joQQ+VQsd/
Lc/+lLcy+0CXiglvrQwyYfZTzwgRwwz55WVKA26YEdYt6KPnmpjOyoBIqPe8OQtaH7voehtzwv+/
AdZLjiDnWbPP20tP5UcjZZxeveuPNec6x7SrtlvibKF/eQKfNNR177VolpCekce0VwioZY3puwDw
I7CIH7V4VEM9t4lc9AOzrj/4Np5CoD7TDYeXODE8j2Lmb8w/5uo8v/Vh85huEVUq7JNAnbVEURZb
HalmsUbfrbB4qcVUbSt4rc6yqC5iUOsVVNAIhScj0vs8IO/MyfdDbztX+/R5RD7c2Bc1FuouVX8W
TzqC59o3lhRynZGSMJdwkje8NaCjqR3dI++nGamnBN9562rDyfiFg6iZYT+z/oJkeiY9yJB9w5qc
Z1qOe+E5cWJyP8SG7oXHRMMncqnrXykK3PrGBFoLjClQuV/ZEZblgioRs0fvLbprOtV8tR0Fy8Zi
6G3na3hRUoHAE4NCQkD0qZNE4D0CoAgdiXKwbmIxhEtNQ/ugQNYtR2L2Xsq4au8NyLB7UUg7+XtM
E23riLtm0IbIMVdA3ibsfFyROPqMvpzkPIUKAFXjUcdUh/ROkg2N658E/tqjT6lRGvdHjfDiPn+5
KYizDWr7QmEeH4vUXDI86pft3LGwlmmGoyDY+kOWrJo7+GRs8sR7s8fzhjsp5WETD9IKPNJerUF1
1vTS3p65xTaNNSpFJPu/PVC2GPoIMbaCNaXi6xLTD50/U+LnE2fW0XLtQzcuPCunOvgrwgea9bKa
zBqNrS/20D2RkXlwbYsf7wO/BV65aOBHRSgYmvmfDd6OmrcOPiKUohxqtGip6MaO7PNSg3CL2gN/
nnDUNDByVx1QTz24P2EWv8D6F5dFrX1aa1WPu55IBmV4tPPtQC2rPBYvPPuSjVJo2aQ3Xk93FPSI
bWh5l4bX31InvO1t24mER/+2F5GQ9HBp2D/2G2i6yLaBhQtB44Gz1NPMqrMbTUARitbO99mER+RF
GKEpDR3QcIGGkHQ4WB1vpWqbdvwX/wCQpkFmTkZlTVKQ2LxOo9IqaDDD5GMu2fXn8lwSLPad/A9h
ZohIBA0wOxxl3i0pxLZgtKMSyVhMITCWVxGL8hwLW9aEB4Ndrsuw+cFOfBOUt7zyHPQIojNUdCeY
/Ku/I+k88C6aD2MqyFehkU+eY26MwNt5C1cANx1at1Jl7EZhoJiSBcsQJpb1RinbMLyL3vwyiZN8
x8Q1iEGVlCHfD9/5CNV7aVtkJpWc4xrjaSQibX7eKD5TZqfavnDTkJFaJZ/wF0WfLhyncxFMMEn+
qV0PqYVCOM6A817hV4pfYWWmgl40hCQzt+ARzZoPauqNXrMFV2nP7ojSLgsWMktoGiewpIK5XGlP
GGs40l/zZM2SM06yhkZHbLaZnXxrFHuov84XFWlwyLVSCRkKwrRNVRMHj60nMlWekSzuB4q0mQEm
eV5wT3bO5dVQDHsZ6GDxUwdJmJ4QG/gsM8nm7VBNmO9c6qzpowI4JOkWpNvSlMqCmvmAYbehlRdi
9Y4WuJf1SYZXeVk4gJK7WBQhQBwwUVheqkiX4SlMVKjdsKkF7+arKxduaT5BkhbUKoYIJr4pZLUL
2uwcRJNpcuRgyaa+PHgyoLRTdjAiQiOvt0Mi/5aG2l/1jGVQNAjZm0dwsLnmlHpOY+aDYHR/I5Mq
bYS0f47HPl3SP8nTIDXK6iKBao6ibOsg9zI781btW9gfsd4FMAZYyhUaYExBRnLIQMN/I/697+Zf
SaBQbpSU4P8Be653LbNodGvKhJBN6nEv1vGQ2XGwts14Op4GfKWEWEkJSv6EOfdN+rIsHdxd9qXV
ri5yQfsSmaElumTFwW0GfMCba86TWP7JLXUlg9fSwZcQITIcWXd3XOwLPtQyFY3eNyeReFvraAeV
F82Btnt8R3UJWfXN1CRpvpye6+DegEIjFzjD5HPQXVc6bQSqwWtueck3lND0Axj3RxYp1APM84AN
FbSE2a46njD6Zqc8XyvODirbdW36yo2ixH5YI7JQbggTdj81FY87Sb+138PADwk3qnekdYwob6as
rKeNP/3Bfc8Q+/i6aukCMgpN7JL1xvpe9fM+fBI2kCDgg7hAOHy3dyQWFhDMvOVKcXon7hf2eyjd
BAfWW1BbqpfOvY/1HxbMFxHyTbNO7EXi4Dhop7ux8tqQzBxIxn/J38ym0nYzYMYYXb/xAwV9StTW
r9iB7uOwbSGXZpVVfB/ijYckoQCo2HCulXFDOdnfz/wyXtJEueKeLUrCYYLXLVQoBmKQ3WeRMdRV
cXdIeGICpbbWrIE65fN5CdIXDf28JpQtCyJIWLoMJWQyxiinU0SCuXWO1Ya6XJagKg2oyMRUMHd7
khSwMLzVmKmYJPJ9usRm0xYjKk+LieEpmhcLbS4VnclV4mi1hJVmRyKW+7VUGgjQLtNgC5qq10pG
nru4fKOHUu3MlIhRcpfPKSUgwiaIu/Ym7vpSA41IohIhHIA3qpdttMXZRa2m00bfWntXBNIeVIcz
9bQAWuNjmmPmwBvQgsZHZKoh7nGyGfJ7y14F6V/MIQBGMYBrD6342/yK8pM3UxesaPj/nng3aAaf
Uz5fdcGJqxcUxkyjT5noJChmCeRN3WwbQfDHE1bHg7u8iNbDL/GH1AlYxQzHD2yy7QxIwjPZIvLK
XZE1/mD9H8c5waF6eKTXxRboc0/HbM0ksYeNWkBxcQHESYXYPYHx8YBLsX8nyKXFXhgcrRPyg+W9
pLMqzA4TRcUPsezviYCUVXTGGLj7TY4NkxPc3ya0bpK7jd2r0FmhvS9h923YLPdxLDwqrMWa6pra
JaNgqDTCMaSI7UO0Tz8owOaXGV3AuwJpzFaHCyjtz1wqEBAYaMZjjDxoH0tXP7kPFV+p1QkLfPST
FMTyoPCZZFFv15CO4lj6qDciOBLCSMOOtNfOT5RzrHIovQVXB6AUHsK4TmRM2S+fnQvHMONZ6crd
WIDIEPxU3Bt++FuJg9jl5yPLOnqDdjV+2K7jySV6boEzMheSdkbl4/aVCRWnwTxQuU2y/0+yi6mK
w683BgoViYTKzyvl3iENU+gGPaQjy3shXDWMNr8VH7nUOwD6hlM6lBXEZfz+Cm6BnycgS/tgVn2v
mAyYiWiNmXbMnQ9rp8ux3nGOjVq1JWSyhu919WiJq7WY+wy/bcr9bZRYAYzMTFJifaGDehvhlmUE
LCuiCyFcYNJ2KiujVv062of+dK53Z3KH6hINDoZbcTtveXq46Znldw80zmrjBmSgBMDRRiqkmhWx
HcX6lsxaHfP9cOqNv+uMzLLFpu1PNm7vfIjDKG3fHLsvEpZ1C/nLpHkm6ykiWvRuvA8zkPtd3OmH
0ba4dBN78vR98I4cldQ2rwR7t58FpgBPLVuSqbdfXxGl9q3gHtGTiyUd5ETKrz1Cy2m5Yb69NlDO
sm+CFo8NTLd5hwqlb0URKhvdUPpiK6daDebgXVPRdVBpBBXXzYz/NPdlSfxdY/t8AG3WAgzOn6AZ
rLMZzmqqKSwU1nqucmYYf8GIcT3Z52ZV/Yml7qaVLtHeG0JLw4JnryO6hRx9tBZkKU1A60YilELx
k20VtXreY936IuI1pPo6MzYiNH9khl033t303Tmu00J4H4B+K9dZgmNoNRhwsVnd+f/qqKqpkpd7
GbipO1Ex7Au45YffnfCGAD6JTDvFHez2LS0wB8CuHKFuOK12bcpP/eTvK6/Y/k7eJWWR9aBfysQq
dx8uojuOnSjpvipDv3sPvn1W4lizLgJ4059//quXBPm5Ujj6BJ37fU01+VBYT6gJnM5dDsH3BY6v
HQhqX7+NmdpQhMgN/eV5fn6VzyvDDI2Bi58XB08z7QJZ8yafRCQnlTKVsJOU8PHIKQ1zkfm4t2bW
QwB4jsFgMGVd8IdFPICmp0AQxOqjf+0oYzfpjQu6WvhVO8RGNTQNA4GmN84Nzn/kECW0e1RsWWTq
0ECPMfrdXLxonRRuAobtoyg8bE5OGDZWnbapbRRFDGgEqh/dDBHlLw2gTHwJPfxDuh/4XJsukF6L
64eLmY4dho7N2NeH6jQ6qzFpwErGP5c8UY/+AKsHNmoeHVAddHwgzHhlp5sJXjNglvLyuBlhR5sr
XaA32oymjvXkBx54Wz3BS+MWK2Aaqtes/nC93rnzx3xY1+Df85O3CFVQoMH3pqbYx9Qpmdw6d1xI
6pxe9a7YwPwzXsRhYOwHRcSIlRJbQnCjRDFWn2QVbCLl3Z+mqkeqyzN0yifRi5Pv/IzJqCb2iV3c
91miouIQyM9tcHs2FDhaG3+NmfoHp+Ov6F+vfKoNdr5CzBd3qoiG4i2UIBgTKE+iipMYrn4LX6J0
F5IVaK+K+7g3tXaSXa2hljS6ifCxnwEQqPYVFhJB+y41Y3wqGQt9JNL5WEp3EqwO63ChXUEcVmWf
/8H0lbBFnrFvg/rl3Ke+n30FOg8oXYbYFxY1Fot9E4b08oqHvcFKVZXGiyw524sPKBvD812sU+48
U0wVJlHIBrYXwzLFCO1pPtykfsiSwn+Rd/wC4XEbkRCpTNFQqnpNVuSMeTCGPD82FsDt4b23Pe1q
hFpNlVCAX2yFakpI/oD0tytxVvngrAiS8dzkX6A4IKWkY/tw35b3qPtBEUggBv0VK3U73QR+f6yh
7o4L7D3qskc7q5Be2imtyX+icE2+61qRMsvEf4iQNW/y2H36b/55ReZCscZrXKVz9/VDhD2yjua2
l+5ScG8xjt2Wy78hayZBfPh9k4uEL2bggNdB59XY5ki+rkip50PRKSh9TxszOdwilijeKdiw70+k
DiqOzEoL/BVLhEOp7P9sNF+MxA90Vra3ToKGtn3VKl8t4RBIOixppx++kJwhjzcJIwBsXwSOc0zP
1Z02vQKIlACVth1V/3lg/18455SGM1ELGl5owtD8kbAorFsQyF7woTAWvGc6HPV2/dIv5ksX+gFo
d0OdjRLvGPxjdFzldpbGj+CU31VuCzFq5e72FHXcdBbg1Ox+OGLygXVX1nF2Jp16oTxihGNJccbs
tvCeY4tNSoijArJn7SUQi8Y0S9wrQGgEKmucJu3vgfl4BuNPwxDgsIoeK1koawl27+7BXADavnCt
LI/p6fhXePgNGY428tpGl0d1H0kzYB1SG4SGng51KodpbssrAzAxZ/C1L1hYyYtP0uIQPookGvJ3
SFIQHX5gNy8KE6GZEj+9+N6mTNH7D+WRP/1d0ZDfb0eAylE3B6x8QqLoHoTSbzQG4Zk4fMLhwNK4
0eug+BC10Uj+yDj85AAKHM7QiSiytLuqoIeqtOB6Ykx2zI7oD1nyT35ggI/zYdePjjlVh2gz/e/Q
kLzf/rpsxQCzC2NM0DQpKpXjKhxozN3KxVzTGP89AT/WmhkK4xy/23Lo2f2Xk2C3kzW9/VKDOTe4
pqmR/mXqEuXmYZ0OuiPOUlatYTaZfffqOI3YSGV5b9urMTlZ4sU6fN1P7OGRHvHkaRyre1d0oqoA
UVT8zVhTun2Edo9/FHCOrVQYXdM4aVT8+AIxzkWhluMeAztsCQWX7DtlXoSsiQfra/5HdEL6h8N1
Xqrp9P25YykuHuFXHMugEEVy63sSwZmYityX5s3aeEx47m3u12mrkNGg422Wu4OKOq1f++m92GY8
xrr+pKPpKH3gWoOpIQdWFHJYkSt8nBhb9DyF9v4KFnXT94597FuIKUqp0Xtpe/a73zaqW1GMB7W+
O4JbAmxoJkftX/f3IYdrLnN8u8+hcmHmdspaDbcpTPr3AStYayNL4FR+rJkRK8wRRXX0wvpxQ4Iy
ocUFjH0tWdpevJWR5rR78rqMzphsQ7JZ/nGPEXLnyapf9gCFUQvGezRKnIWgCzq9xa7Hl7k0v6rl
YzYIDWHHUDxHGhsuwsdOJPnvWhjE7rM9ZswCtrXwezFVY1pesDl7af8lBCvT2DSWzbZ73htObuct
taxi1qcMBD6Q4/X0iK4rogCTEuvKxYwhviXLpm35wk3XrfIEZ617LqgESO5hhgvrHvGOd74g/s3U
Hi+p6byYKvQAgdW0U3cdvvt9N0T13GjMc+/ZfAf6+yUnjfNrPC8uEundXwJenupb/eYAXdP04RJu
1vhymnAqP8M/E2eqjM0+mosiMgNh/oi5YgcvRQh0IK/JGPGSZYu7siVuhJ0T4SmjLW45cQXQiMf8
I6UIg23ASgdipbRszWXlifYxn9IotMojnotrsJ5aTZvOWDpAdHy4rJzUaNufAWuheEnKJtwDkbKA
E2xVzP4gszyLplK3bniAbj8CxiDmGsMI+BnFE5reEn7OhTOTB6EVWpI5tKSySatZUTSCMkjzbga0
BTDM0UXsKMX/UdPgQmZYz7XUsHGVobkW40ma8O3q8I8dCTeOcJAPUGslW8YA5DI3EAeoGGGGsmuJ
7aw5n7c=
`protect end_protected
